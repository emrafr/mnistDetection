library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std;
entity rom_weights is
    port(
        clk : in std_logic;
        romAddress : in std_logic_vector(10 downto 0);
        weights1 : out std_logic_vector(31 downto 0);
        weights2 : out std_logic_vector(31 downto 0);
        weights3 : out std_logic_vector(31 downto 0);
        weights4 : out std_logic_vector(31 downto 0);
        weights5 : out std_logic_vector(31 downto 0);
        weights6 : out std_logic_vector(31 downto 0);
        weights7 : out std_logic_vector(31 downto 0);
        weights8 : out std_logic_vector(31 downto 0);
        weights9 : out std_logic_vector(31 downto 0);
        weights10 : out std_logic_vector(31 downto 0)
    );
end rom_weights;

architecture behavioral of rom_weights is
signal data1, data2, data3, data4, data5, data6, data7, data8, data9, data10  : std_logic_vector(31 downto 0);
type mem is array (0 to 13549) of std_logic_vector(31 downto 0); --change dimension here to 13549 for 10 weights files
constant my_rom : mem := (
0 => "00000000000000010000001000000010",
1 => "00000001111110110000010000000000",
2 => "00000110000000001111111100000010",
3 => "11111111111111011111110111111101",
4 => "00000100000001100000010100001000",
5 => "00000100000000100000000111111110",
6 => "11111100000000110000000111111101",
7 => "00000101000000010000001011111101",
8 => "11111101000000111111111000000000",
9 => "00000010111111010000010111111101",
10 => "11110010111111011111111111111001",
11 => "11111101000000011111101000000011",
12 => "11111101000010111111110111110111",
13 => "11110101111111011111111011111110",
14 => "00000000000000011111011000000100",
15 => "00000010111111100000000100000010",
16 => "11110000111101011110101111110100",
17 => "00001001111110110000100111111000",
18 => "11101100111110101111111011111001",
19 => "11111110111011011111100100000011",
20 => "11110010111011111111001111110111",
21 => "11100110000000111110101100000001",
22 => "11111001111111001110101100000000",
23 => "11111001111101001111110000000100",
24 => "00000011111100001110110111101111",
25 => "00000111111101110000100111110100",
26 => "11110100111101000000000111110101",
27 => "11111101111101011111011100000000",
28 => "00000010000001101111111111111100",
29 => "11101110111011011110111111111110",
30 => "11110000111011011111000100000100",
31 => "11110111111010111110111111111011",
32 => "11101101111000010000100011111010",
33 => "00000101111001100000001111110010",
34 => "11110001111101110000100111110010",
35 => "11111111111001111111011111111111",
36 => "11110001111010110000001011111000",
37 => "11111110111010101111011111111011",
38 => "11100101000000111111011011111111",
39 => "11111010111111001110101100000011",
40 => "11110111111011010000101111111010",
41 => "00001001111001110000110011111000",
42 => "11100110111011110000100011101111",
43 => "11111010111101111111110011111110",
44 => "11110000111010100000000011111001",
45 => "11111001111001001111001011111101",
46 => "11110100111110111111010100000000",
47 => "11110000111111001111111100001001",
48 => "11111011111110110000010111111010",
49 => "00001010111000110000110011111001",
50 => "11101000111010110000101111101101",
51 => "00000111111101101111010100000100",
52 => "11110110110111111111100000000000",
53 => "11111000110111111111110000000011",
54 => "00000101111101111111101100000101",
55 => "11110110111110000000101100010000",
56 => "00001101111100100000001011110001",
57 => "00001011111011100000101011110101",
58 => "11110011111011100000100111110100",
59 => "00000011000000011111101000001110",
60 => "11110100111111001111110011111101",
61 => "11110110111100101111011000001001",
62 => "11110000111100111111011000000000",
63 => "11110100111100111111000100001000",
64 => "11111010111110011111101011110010",
65 => "00001010111101000000111011111000",
66 => "11100111111110000000011011110011",
67 => "00000000111110101111010100000010",
68 => "11110011111101001111011111110110",
69 => "11110001111100001110111000001101",
70 => "11101011111101101111000000000011",
71 => "11110010111011101111101100000101",
72 => "00000000111101001111011111110100",
73 => "11110110111110000000010011110110",
74 => "11111110111101101111111000000010",
75 => "00000000111110111111100011111101",
76 => "11110111111010001110111011110100",
77 => "11101011111101101111100100000001",
78 => "11110001111110101110110000000100",
79 => "11110101111100001111010011111100",
80 => "11111000111101111111100011110001",
81 => "00000010111110110000100111110001",
82 => "11110101111110010000010000000000",
83 => "11111010111110011111001000000000",
84 => "11110000111100101111100111110101",
85 => "11110010111101011111110011111110",
86 => "11110010111101101111000111111110",
87 => "11111010111101111111011011111011",
88 => "11111110111110101111110011110110",
89 => "00000010111110100000001111110111",
90 => "00000100111111011111111000000010",
91 => "00000010111110111111110100000001",
92 => "11111011000000001111111011111101",
93 => "11111101111110101111111100000000",
94 => "11110100111111011111010000000001",
95 => "11111001111101011111010000000000",
96 => "00000010111111001111111000000011",
97 => "00000110111110110000100011111110",
98 => "11111101000000100000001011111011",
99 => "11111101111111100000001111111111",
100 => "11111111111110010000000100000111",
101 => "11111110111111000000000011111110",
102 => "00000001111111101111101111111110",
103 => "11111101000000000000001000000100",
104 => "11111101111111110000001011111101",
105 => "00001010000000100000011100000100",
106 => "11111010000000110000111111111100",
107 => "11111110000000110000010100000010",
108 => "11111111111111100000001111111000",
109 => "00000111000010011111111100000100",
110 => "11111111000001010000011011111110",
111 => "00000001111111111111111000001011",
112 => "11110101111101001111011111101010",
113 => "00000011111001011111111111110111",
114 => "11011001111100000001000011011111",
115 => "11111101111100001111010111111010",
116 => "11110101111110011111001011110011",
117 => "11110011111001001110100011110111",
118 => "11111100111001101110111011111101",
119 => "11110100111001111111101011111101",
120 => "00000010111000011111110011111101",
121 => "00000000111110101111111011110001",
122 => "11110111111100100000000111111000",
123 => "11111011000000101111100000000001",
124 => "11110010111001110000000111111100",
125 => "11110011111100100000011011110101",
126 => "11100110000000101111010000000001",
127 => "11111000000000001110110000000101",
128 => "11111000111010010000010000000110",
129 => "00000110111101100001000011111101",
130 => "11110111111110010000011111111011",
131 => "00000010111110111111110111111101",
132 => "11110101111010111111101100000101",
133 => "11110110111111111111101111110000",
134 => "11110110000001010000000011111111",
135 => "00000001000001011111100000000000",
136 => "11111101110111110000100011111000",
137 => "11111011111111100000010011111101",
138 => "11110110111111000000000111110111",
139 => "00000111000010011111111011110110",
140 => "11111010110110011111110111111110",
141 => "00000001111101100000100011101000",
142 => "11110111111110111111011000000000",
143 => "00000101111101111111110111111001",
144 => "00000000111011111111100111111100",
145 => "11111110000010001111110011111111",
146 => "11111101111111101111111011110011",
147 => "00000010000000101111111000001011",
148 => "11110100111011100000001111110110",
149 => "11110111111111101111110000000000",
150 => "11111010111111101111101011111111",
151 => "00000101111110110000010011101111",
152 => "00001101000000010000100000000000",
153 => "11110110000011110000000111111110",
154 => "00000000000010111111101111111111",
155 => "00000000000100110000001111111100",
156 => "11111101111110100000011000000010",
157 => "00000100111110100000111011110110",
158 => "00000010000010000000100100000100",
159 => "00000101000000111111101111111001",
160 => "00000010111111111111110111111110",
161 => "00000101000001011111111011111111",
162 => "00000010000000000000111111111111",
163 => "11111111000001011111110100000010",
164 => "11110100111111010000010000000011",
165 => "11111010000000010000000100000001",
166 => "11111001000001110000101000000010",
167 => "11111111000001011111111100001000",
168 => "11111011111101001111110000000001",
169 => "00001010000001010000011011111111",
170 => "11111000000001110000110100000000",
171 => "11111111000011010000000011111001",
172 => "11111000110111111111101100000001",
173 => "11111111111011110000100100001100",
174 => "11110000111110100000001000000001",
175 => "00000111111110011111010100001101",
176 => "11111001000001111111101000000001",
177 => "11110110111111100000010111111011",
178 => "11101001000001100000010111110001",
179 => "00001101000001101111110100001011",
180 => "11111110000000000000100011111011",
181 => "00000110111101010000010100000111",
182 => "00000111111111110000111000000101",
183 => "11111110111111001111101100000110",
184 => "11111011111111000000000100000001",
185 => "11100100111110001110111011111101",
186 => "11110111000000011110010011111110",
187 => "11111110111011110000000000000110",
188 => "11111111111011100000000100000001",
189 => "11111101111110011111111111110100",
190 => "11111101111111110000000000000010",
191 => "11111111000000000000011111101110",
192 => "11111100000001011111011111111010",
193 => "00000010111110110000011011111001",
194 => "11100011111110010000100111101110",
195 => "00000101111100101111100111111101",
196 => "11110100000011111111110111101010",
197 => "00000111111110011111011100000111",
198 => "11111001111101110000011000000011",
199 => "11111001111101101111101000000100",
200 => "00000000111000011111101111110110",
201 => "00000101000001010000101011110111",
202 => "11110101111101000000111000000000",
203 => "11111110111110101111100000000100",
204 => "11110110111000111110110100000000",
205 => "11100101111110110000000100001011",
206 => "11110011111111111110010100000000",
207 => "11111010111101011111100000001010",
208 => "11111110111110101111101111111110",
209 => "11110011111110110000010111111110",
210 => "11110001111111001111011011110001",
211 => "11111110000000001111110111111001",
212 => "00000000000000111111111100000010",
213 => "00000001111101111111111011111010",
214 => "11111010000000001111011111111101",
215 => "11111101000000001111111011110111",
216 => "11101111111100111110100111110101",
217 => "11101111111110111111101011110010",
218 => "11111000111011001110001111110011",
219 => "00000100111100101110111011110001",
220 => "11110010111100101111111011111010",
221 => "11100110111110111110111011101010",
222 => "11110110111110011110111011111110",
223 => "11110110111110011110111111110001",
224 => "11110000111001011111011111111100",
225 => "11101000000001000000001100000001",
226 => "11111010111111101110000011111111",
227 => "11111100111101111111101011101101",
228 => "11111101111001111111111100000100",
229 => "11101101111101100000010111100100",
230 => "11111010000000110000010000000000",
231 => "00000000000000001111111111100100",
232 => "00000010111010111111101111111010",
233 => "11101101111100001111111100000001",
234 => "11111010000000001110010111110100",
235 => "11111111000000001111111011110010",
236 => "11110011111001111111111011111111",
237 => "11111111111101001111100111110000",
238 => "11110111111110101110111000000001",
239 => "11110110111101001111010111010111",
240 => "00001010111000110000001100000100",
241 => "11011001000010011110001111111110",
242 => "11111111111111011101101011111100",
243 => "00000100000000100000000111010001",
244 => "11111111110110100000000100000100",
245 => "11111000111110010000110111011011",
246 => "11111100000001000000010011111110",
247 => "11111101111111100000011111011010",
248 => "00000111111100000000011100000010",
249 => "11101111111101111110101100000011",
250 => "11110000111101111110011111111010",
251 => "11111110111111000000011011001010",
252 => "11111001111010111111101011111001",
253 => "11110110111111011111101111011001",
254 => "11111111000010010000100111111011",
255 => "11111010000000000000111111100111",
256 => "11110111111011100000001100000001",
257 => "11111111000001111111111000000001",
258 => "11111100111110011111000111111010",
259 => "00000101111111010000000011110001",
260 => "11111100111100101111111100000001",
261 => "00000000111101111111101011110001",
262 => "11111000111111101111111000000001",
263 => "00000101111111100000001011111010",
264 => "00000001000000001111110100000010",
265 => "11110111000001111111101100000100",
266 => "11110101000001011111110111101111",
267 => "00001010000001011111111011111001",
268 => "11111010111011110000000011101101",
269 => "00000001000000111111110111111001",
270 => "11111111111110100000010000000011",
271 => "00000000111110110000010011111101",
272 => "00000110111110100000010011110011",
273 => "11100100000010011101000100000010",
274 => "00000010000000111110100011111100",
275 => "00010010000000010000110000000110",
276 => "00000111110110111111110111100110",
277 => "00000010000000000000111111110111",
278 => "11111011000011111111111000000101",
279 => "11111101000001100000010111110001",
280 => "11111100000000000000010111111001",
281 => "11110101111111101110111111111011",
282 => "11111110111110111111111000000001",
283 => "11111111111100000000000000001001",
284 => "00000111111011101111111111101011",
285 => "11111011111111000000000111111111",
286 => "11111011111111111111111011111111",
287 => "11111111000001001111101111111010",
288 => "11111101111111100000101111111100",
289 => "11111001000110001110101100000011",
290 => "11101001000010100000001111110100",
291 => "00000110000100110000011000010000",
292 => "00000110111011010000100011101100",
293 => "00000111111110000000110100001011",
294 => "11111111000001010000011000000100",
295 => "00000110000001100000010100001010",
296 => "11111011000101000000001111111111",
297 => "11111000111100011111111111110110",
298 => "11010011111110101111101111101001",
299 => "00000001000001111111110011111011",
300 => "00000010000011010000101011110000",
301 => "00010110111101001111000011110010",
302 => "11111000111101100000101011111111",
303 => "11111100000000011111100111110001",
304 => "11110101111101101111010100000010",
305 => "11011100111011111110000011111000",
306 => "11110001110110011110000111111001",
307 => "00000101111000111111001111111111",
308 => "11110101111010010000100111111111",
309 => "11111110111110101111001111101100",
310 => "00000001111100110000001011111111",
311 => "11111000111100101111101011110000",
312 => "00000011000010001111100111111110",
313 => "00001110111111100000010011111101",
314 => "00001010000001100000001100001000",
315 => "11111101000000001111110100000000",
316 => "11111010000010110000111000001010",
317 => "00010100000001001111111111111101",
318 => "00000000000001000001010100000000",
319 => "00000000111111010000000011111110",
320 => "11110001000000111110111111110011",
321 => "00000110111010010000011111110101",
322 => "00000010111100010000110111110110",
323 => "00000100111010001111000100000001",
324 => "11101010000010011111111111111101",
325 => "00000101111101111101110111110111",
326 => "11110010111010001111010100000100",
327 => "11110001111100011111000111111001",
328 => "00001010111010000000000100000001",
329 => "11101011000001111111110000000100",
330 => "11111010111111011110110100000011",
331 => "11110110111111011111110111110000",
332 => "00001100111010100000000111111101",
333 => "11100100111110100000100111101110",
334 => "00000000000000001111101111111110",
335 => "00000000111111110000001111110000",
336 => "00000000111101111111111000000100",
337 => "11110010000001001110101111111001",
338 => "11111101000000001111010111111110",
339 => "11110100111110110000000011110001",
340 => "11110100111001110000001011111100",
341 => "11110110000001001111001011111011",
342 => "11110100000000111111101100000001",
343 => "00000011111111111111011111101101",
344 => "00000010111110110000000000000100",
345 => "11101110000001101101101100000100",
346 => "11111110000010011101111100000000",
347 => "11111001111111010000010111100101",
348 => "00000111111001001111101111110101",
349 => "00001101111110010000000111110011",
350 => "00000101111111010000001000000001",
351 => "11111111111111110000010011110011",
352 => "00000100000001100000000111111001",
353 => "00000000000010011111111011111111",
354 => "11110011111111101111001111110100",
355 => "00000110000000100000001011100100",
356 => "11111000111111101111000111110100",
357 => "11101101111101011111110111110100",
358 => "11111000111110101111101000000100",
359 => "00000000111101110000001011110111",
360 => "11111111111111100000010111111101",
361 => "11111001000011001111000100000001",
362 => "11110001111111111111110011110100",
363 => "00001001000000110000001011111110",
364 => "00000010111101101111110000000001",
365 => "11111010111100100000010100000000",
366 => "11111110000001000000000000000111",
367 => "00000111111111100000011111111011",
368 => "00001001111101111111101011111001",
369 => "11111111000010001110100100000001",
370 => "11110111111111101111101011111010",
371 => "00100100000010000000001000000010",
372 => "11111011111000110000000111110111",
373 => "00000101111110010000010000000010",
374 => "00000010000001110000010011101110",
375 => "00001000111110010000000000000100",
376 => "00010000000011110000010111111011",
377 => "00000001000111001110110000001110",
378 => "11111000000001100000101111111011",
379 => "00010111000100010000100100011011",
380 => "00000011111101000001001011100001",
381 => "00011000000010100001100100011010",
382 => "00000111000010110000111111011011",
383 => "00001000000001110000010000001111",
384 => "00001000000010100000000011111001",
385 => "11100111000100001100001100000001",
386 => "11111111000001111111011100000100",
387 => "00001001000100110000101000001110",
388 => "00000111111100000000010111011101",
389 => "00001110000000100001010000000111",
390 => "11111100000011000000010011110111",
391 => "00000101000010001111110111110110",
392 => "00001000000010010000101011110111",
393 => "11111101000101001101100000000000",
394 => "11101101000001010000111000000001",
395 => "00000000000000110000101100101000",
396 => "00000010111110100000000111001111",
397 => "00001110111110110001001100011100",
398 => "11111111000010000000011011111011",
399 => "00000110000010000000001100001110",
400 => "00001110000010010000110011110111",
401 => "11111000000100101111001111111010",
402 => "11110011000101100000001011110001",
403 => "11111010000011010000100000001011",
404 => "00010000000000000000001011110001",
405 => "00000110000000010001100100001101",
406 => "00000001000010010000001011111011",
407 => "00001001111111100000000000001011",
408 => "00001010000010010000011111110100",
409 => "11110100111011011111110011110011",
410 => "11110011000011111111101011111101",
411 => "11111111000000011111101000000111",
412 => "00000010000001000000101100000000",
413 => "00001011111101010000100000000001",
414 => "11111100000001011111101000000001",
415 => "11111100111101101111110111111101",
416 => "11111111000010111111111000000001",
417 => "00010111000000000000110011111110",
418 => "00001000000001000001011000001101",
419 => "11111110000000010000000100001011",
420 => "00000011000011100001000100010011",
421 => "00010110000001100000100000001010",
422 => "11111101000000000001110111111110",
423 => "00000000000000010000001100010010",
424 => "11111011000001111111010100000101",
425 => "11111111000001100000100011110011",
426 => "00000011111110011110101011111111",
427 => "00000000111111011111010000000010",
428 => "11110010111111100000010000000100",
429 => "00001010000001101111101000000100",
430 => "11110100000000001111101100000110",
431 => "11110111111111011111011111110001",
432 => "00000001000001100000101100001100",
433 => "11110001000010001111100000000010",
434 => "00001101000011111110110100001101",
435 => "11110011000000110000011011110110",
436 => "00000110000000001111100100000111",
437 => "11110011000010100000011111111000",
438 => "00001000000001010000101111111011",
439 => "00000010000001010000001011101100",
440 => "00000001111011111111110000000001",
441 => "11110001111100011111010011111101",
442 => "11111111000000111110011111111000",
443 => "11110000111110010000011011110010",
444 => "11111011111101001111111111111110",
445 => "11111011111111111111011011110101",
446 => "11110101111111000000001111111101",
447 => "00000110111111010000000111110100",
448 => "11111101000001000000000011110111",
449 => "00000011111111100000111000000001",
450 => "00000011000001111111110111111100",
451 => "11111100000000101111101011111011",
452 => "00000110000010101111010100001000",
453 => "00001001111111011111100100000100",
454 => "00000111111111001111011011111111",
455 => "00000010000000001111111100000001",
456 => "11111101000000101111110100000000",
457 => "11111011111111001111101111111101",
458 => "00000010000010101110111011111101",
459 => "11110001000010011111111011110001",
460 => "11111100000001111110101011111011",
461 => "11111001111110001111100011111011",
462 => "11111011111110100000000000000110",
463 => "11111111111111100000001111111110",
464 => "00001101000011100000000111111110",
465 => "11111100000110001110100000000000",
466 => "11111101000000101111010000000011",
467 => "00000111000011110000100000001000",
468 => "00000010111110001110001011110010",
469 => "11101010111111010000101111111000",
470 => "00001011000001001111011011111001",
471 => "00000100000001010000010111111000",
472 => "00010010000010100000011111110010",
473 => "00000000000101001110011011111001",
474 => "00000001000001001111110100000011",
475 => "00100001000011100000000000001011",
476 => "00001010111101001110000111011111",
477 => "11101111000001000001000100001111",
478 => "00000110000011011110010011101110",
479 => "11111110000010000000010011111100",
480 => "00001001000110000000010011110001",
481 => "11110101000010001110000111111100",
482 => "00000100000001011111110000001011",
483 => "00110000000001010000001000001011",
484 => "00001000111101111111100111001101",
485 => "00010101000010010001100000001100",
486 => "00000101000010101110110111111000",
487 => "11111100000000010000000000001000",
488 => "00001110000110010000110111110001",
489 => "11101101000100011100101111111111",
490 => "00010001000001011111110000010111",
491 => "00001011000010101111111000101000",
492 => "00001111111101011110100011010001",
493 => "00001010000100110001011000010000",
494 => "00010100000011001101110111110000",
495 => "00000011000011000000100100000010",
496 => "00000001000101000000011011111001",
497 => "11101010000100111101100000000101",
498 => "00100100000001101111001100011111",
499 => "00001010111111111111111000011011",
500 => "00000010111111111111000111001101",
501 => "00001101000011010000111011111111",
502 => "11111110000001010000000111101110",
503 => "00000101000010110000001111111010",
504 => "00000001000011010000010011111110",
505 => "11111010111111101111000000000101",
506 => "00011111000001011111101000011100",
507 => "00000011000000011111100000001101",
508 => "00001101000001111111101011100111",
509 => "00001100000011010000110100000110",
510 => "00001110111111100000000111110101",
511 => "00000011000011000000000111110111",
512 => "11110111111111111111110111110100",
513 => "11101101111101001111000111111111",
514 => "00000001111110011110000111111100",
515 => "11111010111110011111101111111100",
516 => "11111100111111111110101100000000",
517 => "11110111111101011111010011110000",
518 => "11111101111110001111001011111110",
519 => "11111110111110101111101011100000",
520 => "00000011000011000000001011111011",
521 => "00010000111111110001001011111111",
522 => "11111101000000110001011100000010",
523 => "00000000000001011111110000001000",
524 => "00000001000011010000011100000101",
525 => "00010110111101010000001100000100",
526 => "00000001111111001111110111111101",
527 => "11111011111111101111110000001011",
528 => "11101110000001101111100100000000",
529 => "00000010111011000000101011111101",
530 => "11111110000000000001000100000100",
531 => "00000001111100111111111100000001",
532 => "11111010000001100000101111111101",
533 => "11111100111111111111100111111011",
534 => "11111110000000000000010000000011",
535 => "11110111111111101111100111111001",
536 => "00001001111111010000011011111111",
537 => "11100010000001111110000011111111",
538 => "00011010000001011110111100010000",
539 => "11110001111111100000010100000001",
540 => "00000110000001101111101000000101",
541 => "11110111000010110000111000001011",
542 => "00001100000011001111011011111011",
543 => "00000011000010010000011011100001",
544 => "11110001000010011111110100000101",
545 => "00000100111000000000110100000001",
546 => "00001110111111001111001100000100",
547 => "11101001111110101111101111100110",
548 => "00000011000110010000011000001111",
549 => "11111010000001001111100011110011",
550 => "00000111000001000000011011111111",
551 => "11111011000000110000000011101011",
552 => "11111110000001110000000100000101",
553 => "11111110111010100000010011111111",
554 => "00010010000001001111001000010010",
555 => "11011100111111011111111011110010",
556 => "00001000000010111111011100011110",
557 => "11101110000010000000010000000011",
558 => "00010000000010100000101111101111",
559 => "11111100000010010000000111111000",
560 => "00000001000011100000010100000000",
561 => "11110111000001001110111000001000",
562 => "11111101111111011110011011111100",
563 => "11111011000001101111110111110011",
564 => "00001011111111101110010100000000",
565 => "11111000111111110000110111110011",
566 => "00010001000000111111110011111100",
567 => "00000000000001000000101111110101",
568 => "00001000001001001111101111110010",
569 => "00000110000010100000010111111110",
570 => "11110000111110000000011011111000",
571 => "00011011000001001111110100011011",
572 => "11111000000100101101010111110011",
573 => "11101101111111010000100100000110",
574 => "00001000111111011101111100000011",
575 => "11110101111111011111111000000011",
576 => "00000100000111101111100111100010",
577 => "11111110000000101111100011111011",
578 => "00001110111110000000110000010111",
579 => "00010110111110101111011000101010",
580 => "11111001000011101100001011011001",
581 => "11011101000001100000101000010101",
582 => "11111010111110111100111000000100",
583 => "11101111111110001111101000000101",
584 => "00000001000001101111101111101100",
585 => "11100111000001101110010111111000",
586 => "00000111111110001111100100010011",
587 => "11111101111111011111101000001100",
588 => "11111110000000001101000111100001",
589 => "11101011000001000001001100000011",
590 => "00000010111111111101110011101010",
591 => "11111010000001011111100011101111",
592 => "00000001000100010000010111111111",
593 => "11110000000010001101111000001010",
594 => "00010101000010011111001000010101",
595 => "00001001000000100000010000011000",
596 => "00001110000000101101111011011101",
597 => "00000110000011110001000100000110",
598 => "00000111000001011110111011101101",
599 => "00000001000001010000010111111010",
600 => "00001000000100000000011111111111",
601 => "11110110000100011110001000000010",
602 => "00100001000001111111001000011100",
603 => "00000001000001110000110000100000",
604 => "00001000000001011110111011001111",
605 => "00001001000100110000101111111110",
606 => "00001010000001101110111111100001",
607 => "00001101000000100000000011110110",
608 => "00000101000101000000101011111101",
609 => "11111010000001111110111100001100",
610 => "00011011000000001111101000011000",
611 => "11111101000001011111100100001000",
612 => "00010101000101011111110011110000",
613 => "00001111000100100001100000001010",
614 => "00001110000011100000010111110110",
615 => "00000100000100000000100000000000",
616 => "11111011000000101111110111110110",
617 => "11110110111100101111110100000100",
618 => "11111000111010011101011111111101",
619 => "00000101111011100000010011111110",
620 => "11111101111111111111110111101100",
621 => "00000101111101111111101111011100",
622 => "11111110111101011111111100000010",
623 => "00000001111110011111101111101000",
624 => "11111000111111001111011111110110",
625 => "11110100111101110000010111111011",
626 => "11101001111101011111101111110011",
627 => "11111101111100111111111000000100",
628 => "11111001111111010000000011111000",
629 => "00000101111101111111010011111101",
630 => "11111001111101100000001000000011",
631 => "11111001111101111111110111110100",
632 => "11110001000010001111110011111000",
633 => "11101101111110001111111111111011",
634 => "00001011111111111111100000001011",
635 => "11111101111110011111111011111100",
636 => "11110111000001111111011000001000",
637 => "11110011000000011111111100000110",
638 => "00000111000001001110101100000010",
639 => "00000000000000101111110111101100",
640 => "00000001000110010000001100000101",
641 => "11100000111111111110101100000111",
642 => "00011110111111011110110000010010",
643 => "11100100000001100000010111111011",
644 => "00000100000101101110101100000000",
645 => "11110100000101000000010011111110",
646 => "00010001000010001111011011110111",
647 => "00000011000011010000100011100001",
648 => "00000100000101010000100100001100",
649 => "11101101000010001111011100001010",
650 => "00010010000010101101110000010110",
651 => "11010100000001000000100011010000",
652 => "00010111000111001110011000010001",
653 => "11110111000010000001011111101000",
654 => "00001000000101010000001011101111",
655 => "00000110000010000000111011001010",
656 => "00000000000101011111111100000101",
657 => "11111101111101101111110000001011",
658 => "00011000000001101110010100010101",
659 => "11100100111111101111101111011011",
660 => "00001101000011001110010000000101",
661 => "11110000000001111111101111110010",
662 => "00011000111111110000110011100101",
663 => "00000001000001100000011111101111",
664 => "00000100001010100000000011111001",
665 => "11110100000000101111100011111110",
666 => "00000100111111101110010000000111",
667 => "11111000111101111111111011100101",
668 => "00000100000100101100011111101000",
669 => "00000010000000100000110111101100",
670 => "00001110000000101110010011111010",
671 => "11111101000000000000001111110101",
672 => "11111011001011111110110111100101",
673 => "11110100111100111111101011110001",
674 => "11101101111001101110101111110101",
675 => "00011111111010011110110111111011",
676 => "11111011000110001100110011101011",
677 => "11110101111011011111101111110001",
678 => "00000001111100011100111100001010",
679 => "11101111111101011111011111100100",
680 => "11101110000011011110011011100100",
681 => "11100111111100111111000111101100",
682 => "00010011111011101111001100011101",
683 => "00101100111011101110100100011010",
684 => "11101010000000101101010111101011",
685 => "11011111000000001111010100000100",
686 => "11110010111001101101100000010001",
687 => "11100110111101101110101011101101",
688 => "11110010111111001111101011111010",
689 => "11110000111110111110100111111111",
690 => "00010111111110001111101100100011",
691 => "00000101111101111111110100100010",
692 => "00000101111110001100110000000000",
693 => "11011101000011001111111000000110",
694 => "00000011111110111110000111111101",
695 => "11111011000001111111110111111110",
696 => "11111011000001010000100000000001",
697 => "11111111111111101111100011111111",
698 => "00001101111111111111011000001010",
699 => "00001001000000010000000100011111",
700 => "11111111000010001110001011111011",
701 => "11110100000000110000010000000000",
702 => "11111110000001111110110111110101",
703 => "00001000000001011111111000000010",
704 => "00001001000100000000100100000001",
705 => "11111101000010001111000100000001",
706 => "00011110000000101111100100100100",
707 => "11101010000010100000010000010110",
708 => "00001001000100001110011100000111",
709 => "11110100000010010000111100000000",
710 => "00001101000010101110111111101110",
711 => "00000100000010100000011011111001",
712 => "00000111000100110000101100000100",
713 => "11111010000101001111011000001001",
714 => "00011010111110111111111100010010",
715 => "11101011000011010000101111111101",
716 => "00001010000011111110110111110100",
717 => "00000111000100010001111011110110",
718 => "00000110000101101111001111111001",
719 => "00001001000001010000001100000010",
720 => "11111101000011000000010111110111",
721 => "11101011111101001110011011111111",
722 => "11101010111110011101111011110011",
723 => "11111011111010100000001011111100",
724 => "00000010000010010000000011111000",
725 => "00000100111110101111011111100100",
726 => "00000010111101110000000011111011",
727 => "00001001111110100000010011101010",
728 => "11110011111111111111110011110011",
729 => "11011111111010110000001111110101",
730 => "11110011111111001110001011110000",
731 => "11111101111101011111011111110101",
732 => "11111000111111110000001011111011",
733 => "00000001111100001111010111101001",
734 => "11111110111011111111111011111110",
735 => "11110111111100001111001111100110",
736 => "11110010000010011111111100001110",
737 => "11101111000000001111110100000000",
738 => "00001010111111101111010100001101",
739 => "11110111111111011111111000000100",
740 => "00000001000000001111100100000111",
741 => "11111110000000100000001000000010",
742 => "00000011000010000001001111111100",
743 => "11111110000010000000001011110000",
744 => "00000011000101010000011000000111",
745 => "11110110000000101111000100001111",
746 => "00010110000001011111110000011011",
747 => "11100111000000100000000111111111",
748 => "00000010000111111110010000000000",
749 => "11110000000100100000010100001000",
750 => "00000100000010100000010011110011",
751 => "00000100000011100000000111110011",
752 => "00001001000110110000101000000101",
753 => "11110010000010111110001100001001",
754 => "00010111000011101110001100011000",
755 => "11100000000001010000001111101010",
756 => "00011011000011111101110111110000",
757 => "11111000000010110001100111110101",
758 => "00010010000011001111000111100101",
759 => "00001000000010100000110111100000",
760 => "11111111000110010000011111111101",
761 => "11101011111110011111101000000100",
762 => "00001010111111111110000100010001",
763 => "11011111000001000000100011100101",
764 => "00000111000011101101001000000100",
765 => "11110001000010101111100111101111",
766 => "00010101000000101110100111011111",
767 => "00000111000001000000011111100011",
768 => "11111011001000100000001011111101",
769 => "11101110111100111111110011111110",
770 => "00000111111111011110011000000011",
771 => "11110100111001111111110100001000",
772 => "00001001000110001110010111111101",
773 => "00000011000000001111011111101011",
774 => "00001111111101111110111011111011",
775 => "11111011111111010000010011110101",
776 => "11111010001000111110110111110000",
777 => "11101000111011101111010011110001",
778 => "11110011111100001110011111111110",
779 => "00001000111001011110100000000101",
780 => "11101011000110101110111000000000",
781 => "11111110111100101111100111101111",
782 => "11110001111110011111001100000111",
783 => "11100110111101111110100111101010",
784 => "11100100111100001110100011111101",
785 => "11010000111101011110000011110101",
786 => "00010001111111001100101100010001",
787 => "00010101111010001110101111111011",
788 => "11110010111010110000000100010110",
789 => "11101011111111011111110011100100",
790 => "11110111111110010000010000001101",
791 => "11110101111110011111001111010011",
792 => "11110001111101001111001100000110",
793 => "11101010111010101110101000000100",
794 => "00010010000000101110001100010001",
795 => "00000101111100111111011100000101",
796 => "11111101111101111110001111110101",
797 => "11011100000011001111010011101100",
798 => "11111111111101001111111100001110",
799 => "11110110000010001111010111100111",
800 => "11111100000000010000001111111100",
801 => "00000010111110110000000111111110",
802 => "00010001000001001111111000000111",
803 => "11110011000000100000001000011000",
804 => "00000110000001111110101000000111",
805 => "11110001000000110000000000000011",
806 => "00000100111110111110110111111100",
807 => "00000100111111110000000011111110",
808 => "00001011000001110000011111111100",
809 => "00001000000001000000010000000011",
810 => "00000101000000110000001000001001",
811 => "11100111000001000000010100000001",
812 => "00000011000100001110001000001110",
813 => "11101010000001100001001000000100",
814 => "11111111000100101111010011111010",
815 => "00000100000001000000001011111111",
816 => "00001101000101010000101111111010",
817 => "00000110000001100000101000001011",
818 => "11110011000001101111111011110101",
819 => "11111010000000110000100111101101",
820 => "00001011000011101110011000000001",
821 => "00000000111111110001000111111101",
822 => "00001011000001111111000111111001",
823 => "00001001000001100000001100001010",
824 => "11111100000100000000000111101111",
825 => "11110110000001111111110011111001",
826 => "11111001111010101111001011111110",
827 => "11111110111110000000001111111100",
828 => "11111011000011001111010011101111",
829 => "00000000111110110000001011111000",
830 => "11111110000001001110100100000010",
831 => "11111111111111001111110100000100",
832 => "11110100000001001111101111110010",
833 => "11110110111100110000101011111001",
834 => "11110001111101111111000111110011",
835 => "11111111111101111111100111110111",
836 => "11111101000000110000000111111101",
837 => "00000110111101011111000011111001",
838 => "00000000111101100000010111111101",
839 => "11111001111100011111100111111001",
840 => "11111110000011100000010000000001",
841 => "11111111000001110000010100000111",
842 => "00000001000010011111100100001010",
843 => "11111000000010000000000000000011",
844 => "00001000000100011111000000000011",
845 => "11101101000000110000101000000011",
846 => "00000011000000100001001111111001",
847 => "00000010000000100000011000000100",
848 => "00000110000010110000100100000001",
849 => "11111101000011001111110100001011",
850 => "00000111000001111111101100001101",
851 => "11111100000010100000011011111110",
852 => "11111110000001011101011111101001",
853 => "11110111000010001111101100000100",
854 => "11111100000000100000010011110111",
855 => "00001000000010100000011111111110",
856 => "00001110000100100000111011111100",
857 => "11110110000100011110001100001110",
858 => "00001100000010001111001000001101",
859 => "11101110000001010000111100000010",
860 => "00001110000011011110000011011110",
861 => "11111010000010110001000011111001",
862 => "00001100000101111111101111010111",
863 => "00001000000011000000010111110111",
864 => "00000001000101101111110000000100",
865 => "00000001000001001110100000000101",
866 => "00001111000010111111010000001000",
867 => "11100000000000111111111100000011",
868 => "00001000000100101110101111101111",
869 => "11111110000010010000001011110111",
870 => "00001001111111101111101111100100",
871 => "00000010000000110000011111110010",
872 => "11111011001010011111110111110111",
873 => "11110010111110001111110111110110",
874 => "00001101111111011101101100000101",
875 => "11111001111110001111100011101101",
876 => "00000101001000011111011100000101",
877 => "00001001111111011111110111011111",
878 => "00011000111110011111000111110100",
879 => "11111110111110001111110011101100",
880 => "11110001000100101110110000000011",
881 => "11100011111010101111010111110011",
882 => "00010000111110111110010000010010",
883 => "00000101110111011110101011111111",
884 => "11100111000001111111110100001101",
885 => "11111111111111111110110011101011",
886 => "11110001111101010000101100001001",
887 => "11110000111110101111011111101001",
888 => "11100100111101011111000011111110",
889 => "00000001110110110000011111111111",
890 => "00010000111111101110110000001000",
891 => "00000110111100011111000011101011",
892 => "11110000111110111111110000010011",
893 => "11100100111110101110000111101001",
894 => "11111110111100100000000100000110",
895 => "11110111111110111111110011110101",
896 => "11111001000000001111100100000100",
897 => "00000101111101010001011000000101",
898 => "00000011111111010000001100001010",
899 => "11110011000000011111000111110110",
900 => "11111100000001111111111100010000",
901 => "11110110111111011111011111111101",
902 => "11111011111100010000011100000001",
903 => "11110111111110011111101100000011",
904 => "11111011111111110000000000000110",
905 => "00000111111011110000000100000110",
906 => "00010101111111001111110000011001",
907 => "11111011111101101111110011110111",
908 => "11111001000000101110110000011000",
909 => "11101011000010011111100011111110",
910 => "11111111000001101111100100000100",
911 => "11111100000001101111111100000000",
912 => "00000011000000001111101100000000",
913 => "00000101111111100000010000000011",
914 => "00001010000000000000000000001101",
915 => "11110001111111100000011111111001",
916 => "11111100000000111110010100001111",
917 => "11101001000000100000000000000110",
918 => "11111100111111101110111100000001",
919 => "00001010000001110000010011111110",
920 => "00001000000001000000100011111101",
921 => "00000111000011100000010000000110",
922 => "11111111111110111111110011111001",
923 => "11110000000001100000101111111011",
924 => "00001101000010111101011111111011",
925 => "00000010000000010000100100000000",
926 => "00001101000001011101111100000001",
927 => "00000111000000100000001000000100",
928 => "11110011000001001111001111101011",
929 => "11110110111100001111101111111010",
930 => "00001000111001001111010111111111",
931 => "00000000111100001111100100000100",
932 => "11110111000001011111010011111000",
933 => "00000111000001001110110011110000",
934 => "11110111111001111111000000000100",
935 => "11111001111101011111110111110110",
936 => "00000000000010001111011111111001",
937 => "11110010111110010000011111110110",
938 => "11111111111110011110101011111000",
939 => "00000010000000001111110011110111",
940 => "11111000000001110000010100000110",
941 => "00001101111111111111110011111111",
942 => "00000010111110011111110100000000",
943 => "11111011111111001111010111110100",
944 => "00000101000110000000011111111011",
945 => "11111110000010101111100100000010",
946 => "11111100000001101111110111111110",
947 => "00000001000010010000100000001010",
948 => "00010011000000011110100111111001",
949 => "11111011000000000000101000000111",
950 => "11111111111111011111110011111001",
951 => "00000100000000010000101111111101",
952 => "00000010000010010000010100000000",
953 => "11110000000000111111010000000011",
954 => "00000001000000111111001111111101",
955 => "11111101000010010000000100000000",
956 => "11111111111110101101101011100010",
957 => "11111000000001010000000100000001",
958 => "11111111111111111111101111111101",
959 => "00000001000001010000011011111011",
960 => "11111101000011000000110011110100",
961 => "11111111111111111111011100000011",
962 => "11111001000000111111110111111110",
963 => "11110000000001010000011000001011",
964 => "00000100000100001101001011010110",
965 => "11110001111111100000000000000000",
966 => "00010000000001011110000111111010",
967 => "00001000000001100000100100000001",
968 => "00001011000110110000111011111110",
969 => "00000010000011011110111111111111",
970 => "00010001000000010000101000001000",
971 => "00000101000000011111111100011001",
972 => "00010001001000111111010011111000",
973 => "00000011000011000001011100001010",
974 => "00010011000011101111011011011110",
975 => "00000010000010010000001100010001",
976 => "00000101001000001111101100001000",
977 => "11111100111111111111110100000110",
978 => "00011010000000011111111000010110",
979 => "11101001000000000000010100001111",
980 => "00000100000010110000000111111101",
981 => "00000011000100000000111000000011",
982 => "00001010000100001111111111101001",
983 => "00000111000000011111111100000100",
984 => "11110010000010111111001100000011",
985 => "00000010111011000000111100000011",
986 => "00000111111111110000011000000000",
987 => "00001100111110001111111111111111",
988 => "11101101000010100000010111111000",
989 => "11111010000000111110010111110010",
990 => "11101100111110010001001011111111",
991 => "11111011111101111111101011111111",
992 => "11110000111111101110110100000111",
993 => "00000111111001000001110011111110",
994 => "00000101111111000000100000000111",
995 => "11111000111011101111011111110000",
996 => "11110001000010010000101000010001",
997 => "11110110000000111110010111110110",
998 => "00000001111110010000110011111101",
999 => "11111101111110111111101100001011",
1000 => "11111000111011001111101000000010",
1001 => "00000000111011110000011000000011",
1002 => "11111110000000101111110011111111",
1003 => "11111101111100111111101111100010",
1004 => "11110101111110110000000100001100",
1005 => "11101110111111001110000111110011",
1006 => "11110010111011100000100000010011",
1007 => "11111101111101011111101000000010",
1008 => "11110010111101011111011111111111",
1009 => "00001001111100000000100100000010",
1010 => "11111010111111011111110111110111",
1011 => "11111101000000010000000011111110",
1012 => "00000000000000011111001111111010",
1013 => "11101111111101101110000111111101",
1014 => "11111010111100111111101000000001",
1015 => "00000010111110010000000000000111",
1016 => "00000001111101111111111000001100",
1017 => "00001100111111010000111000000101",
1018 => "11111100000001101111111000001011",
1019 => "11110100000010011111111011101101",
1020 => "11110111000000101110010000001010",
1021 => "11100110111111010000000011111100",
1022 => "11110101111101111111110000000110",
1023 => "00000010111111100000010000000110",
1024 => "00000101111110111111110111111011",
1025 => "00001010111100010000011100000111",
1026 => "11101010111011001111101011110111",
1027 => "11111101111110010000100111100010",
1028 => "11110111000001001101110100000001",
1029 => "11100110111101101111011011111100",
1030 => "11111110111111011110111000000100",
1031 => "00000010111100110000011011111001",
1032 => "11111001000000111110111011110101",
1033 => "00000000111110000000101011111011",
1034 => "00001001111001001111100000000011",
1035 => "11111101000000111111101111111100",
1036 => "11110011000000001111100000000101",
1037 => "00000000111110111110110111110111",
1038 => "11101101111111011111010100000101",
1039 => "11111001111110101111011111110100",
1040 => "11111100000000011111111111111100",
1041 => "00000111111101100000000111111010",
1042 => "00000000111101110000100000000100",
1043 => "00000001111111001111111000000000",
1044 => "11111111000011000000000000000001",
1045 => "00000010000000101111111100000110",
1046 => "00000001111110111111111111111110",
1047 => "11111101111111101111011000001011",
1048 => "00000110000000100000000111101011",
1049 => "00000011111101100000110111111110",
1050 => "11111111111101100000001111111101",
1051 => "00000101111111000000010100000011",
1052 => "00000011000000001110101011100010",
1053 => "11101011111101110000000111111110",
1054 => "11111111111100101101101100000011",
1055 => "11110110111111000000001111111011",
1056 => "11111110000000010000011011111101",
1057 => "11111001000000011111100111111101",
1058 => "00001100111111101111101100000010",
1059 => "00000001000000011111111000000101",
1060 => "00000101111100011101010111011010",
1061 => "00000001000011010000001000000010",
1062 => "00000111000000011101110011111101",
1063 => "00000011000001110000010111111100",
1064 => "00001101000011000000111011110011",
1065 => "11111001111111101110111000000100",
1066 => "11110010000001011111110011111010",
1067 => "11110110000000110000100000000001",
1068 => "00000111000011001110000010110001",
1069 => "11111110111110110000101011111101",
1070 => "00001110000000001101111100000010",
1071 => "00000110000001000000000100000000",
1072 => "00000011001001000000100111110111",
1073 => "11111110111111101110001100000001",
1074 => "11111111111110110000000000000001",
1075 => "00100100111110110000010100001011",
1076 => "00001101000010111111011011011001",
1077 => "00001011000010000000100100001010",
1078 => "00000100000001111111000111111110",
1079 => "11111101000001101111110111111110",
1080 => "00001100000010110000011011111011",
1081 => "00000001000010101111001100000011",
1082 => "11101101111111110000011111101111",
1083 => "00110000000000111111110000001110",
1084 => "00000111111101100000010111110001",
1085 => "00001001111110110001010100000101",
1086 => "00000100000010001111101111111001",
1087 => "00000100000001000000010000000011",
1088 => "11111111111010001111010011111101",
1089 => "00000011000011100000010011111101",
1090 => "11100000111110010000110011011001",
1091 => "00100010000010010000000111110100",
1092 => "11110101111001010000101100011011",
1093 => "11110111111100110000010111111110",
1094 => "11101101000010110000010100001110",
1095 => "00000010111111111111110000000110",
1096 => "11111111110111001111101000000110",
1097 => "00000001000001010000001100000001",
1098 => "11100110111111101111100111100001",
1099 => "00010011111111010000010011100101",
1100 => "11110011111011000000011000000101",
1101 => "11011110111110111110100011110001",
1102 => "00000000111111000000101100001000",
1103 => "11111111111110101111111011111111",
1104 => "11111000111010101111111011111100",
1105 => "00000000111100000000010011111111",
1106 => "11010111111100111111011111010000",
1107 => "11111011111110100000010111010101",
1108 => "11101111111110010000001000000101",
1109 => "11011000111010011101110011110010",
1110 => "11110101111110010000000000011001",
1111 => "00000100111011101111110011111000",
1112 => "11110011111011011111101000001011",
1113 => "11111100111100110000011000000011",
1114 => "11100100111010101111011111110001",
1115 => "11110101111101011111010111100000",
1116 => "11110001000000111111101100010010",
1117 => "11001110111100011110001011110011",
1118 => "11111000111011100000111100001000",
1119 => "11110100111110010000001111111101",
1120 => "11111111111000110000000100001000",
1121 => "11111001111110011111111000000000",
1122 => "11101000111110100000000011101010",
1123 => "11111111111100100000000011101101",
1124 => "11111000111101001111100000001000",
1125 => "11000110111011111111000111111001",
1126 => "11110111111101000000011100000000",
1127 => "00000010111110000000000111111001",
1128 => "11111011111100011111011111110101",
1129 => "00000000111011101111110011110101",
1130 => "11101001111100001111011111101011",
1131 => "00000000111111101111100111100001",
1132 => "11101111111110110000010100001001",
1133 => "11100100111010001110011111101100",
1134 => "11110111111011111111110100000001",
1135 => "11111000111010111111110111110101",
1136 => "11101111111011111111010011111111",
1137 => "00000011111101100000011011111111",
1138 => "00001011000000000000000100000001",
1139 => "00000001111011111111001000000011",
1140 => "11110010111100100000101000010010",
1141 => "11101101000010111110010011110101",
1142 => "11110000111010110000001000000001",
1143 => "11111010111111101111010011111001",
1144 => "00000001000000011111110111111011",
1145 => "11101110111111110000000111111000",
1146 => "11110000111110001111000011110010",
1147 => "00000001111110100000000111110101",
1148 => "11111110111111101111110100000100",
1149 => "00000000111100101111100111110001",
1150 => "11111011111110111111110100000100",
1151 => "00000000111110001111111111101000",
1152 => "11111100111110101111101000000100",
1153 => "11111010111111111111000111110100",
1154 => "11111111111100111111001111111110",
1155 => "00000010111110001111101011111100",
1156 => "11111001111110111111111000001101",
1157 => "11111110111111001111111111110011",
1158 => "11110001000001100000011100000111",
1159 => "11110110111111101111011111110110",
1160 => "00000110111010110000110111111100",
1161 => "00001000000001010000010100001010",
1162 => "00000100111111010000110000001010",
1163 => "00000100000000100000011100001110",
1164 => "00000110111010001110001011010011",
1165 => "11111101000000001111110000001010",
1166 => "00000110111111011111101111111101",
1167 => "11111111000001100000010100000101",
1168 => "00010100111100110001011111101000",
1169 => "00000110000011110000001111111001",
1170 => "11101010111111110000111111110011",
1171 => "00001010000010000000111100001110",
1172 => "00001010111110001111001011010100",
1173 => "00001011111101110000110100001110",
1174 => "11111110000011111110001100000001",
1175 => "00000100000010010000000100010000",
1176 => "00001011111111000000010011110000",
1177 => "00000110000010101111111011111100",
1178 => "11011100111110100000101011100100",
1179 => "00010000000010010000000000000010",
1180 => "11111110111110000000010111100001",
1181 => "00011101111111000001110000001011",
1182 => "11101111000011001111111111111110",
1183 => "00000001111110000000011100001001",
1184 => "00010001111101011111000111101110",
1185 => "00001010000100101111111011111100",
1186 => "11011001111110100000011111100001",
1187 => "00001110000010110000100000000101",
1188 => "11111110111111000001000111111001",
1189 => "00001000111101110001101100000101",
1190 => "11101110000100001111001111111100",
1191 => "00001010111110011111101100001011",
1192 => "00000100110011011111010111111011",
1193 => "00001011000010110000100000000001",
1194 => "10101100000001110000111010110010",
1195 => "00000100000010000000011100000001",
1196 => "11110110111011100010111111111101",
1197 => "00000001111000000000001100001001",
1198 => "11100100000000010000111011111111",
1199 => "00000111111011110000001000001011",
1200 => "00001001110100010000100011111011",
1201 => "00000110000010110000011011111101",
1202 => "10111000111111010000011010110110",
1203 => "00000010000000000000010111110000",
1204 => "11101100111010010001111111110001",
1205 => "11010100110110111111010100001011",
1206 => "11101110000010010001100000000000",
1207 => "00001011111101100000000100001010",
1208 => "00001000111011000000000111110111",
1209 => "00001000000010100000111011111011",
1210 => "10111101000010100000100111000011",
1211 => "11101111000011010000010011110001",
1212 => "11110110111111000010010100001100",
1213 => "11010100110111101111110000000111",
1214 => "11111000000000110001000000000100",
1215 => "00000010111111010000101100010000",
1216 => "00000010111010011111111011111000",
1217 => "11111010111101000000001011111100",
1218 => "11001011111110111111110011010100",
1219 => "11111101111110001111101011101010",
1220 => "11101000111111100000101100001001",
1221 => "11010011111000011110101011111010",
1222 => "11100101111101000000101000000011",
1223 => "11110010111101101111101111111001",
1224 => "11110100110110001111110011110010",
1225 => "11110111111011101111110011110110",
1226 => "11100001111110011111100111100100",
1227 => "11111111111101101111100111110011",
1228 => "11101101111011011111010111111101",
1229 => "11001010111001101111001111111010",
1230 => "11101011111100011110101000000000",
1231 => "11110111111110001111111111111111",
1232 => "11111010111100101110101111110110",
1233 => "11110011111011011111011111101101",
1234 => "11110000111011101111011111110011",
1235 => "11111010111101001111101111100111",
1236 => "11110010111101100000000000001101",
1237 => "11100001111100111111000111110000",
1238 => "11100111111011111111010011111111",
1239 => "11110111111011011111101011101110",
1240 => "11111001111011001111110100000011",
1241 => "11101001111101001110111000000000",
1242 => "00000000111100001110101100000001",
1243 => "00000100111101001111101000000100",
1244 => "11111100111001110000001111101110",
1245 => "11101100111111011111001111101101",
1246 => "11111000111011001111111000000100",
1247 => "11111011000000001111101111110101",
1248 => "11111001111111101111101100000001",
1249 => "11110111000000010000001111111101",
1250 => "11111010000001011111001011111000",
1251 => "00000001000000001111110000000010",
1252 => "11111100000001001111111100000010",
1253 => "00000111111111001111111011111010",
1254 => "11111010111111000000011000000100",
1255 => "00000011000000001111111011111100",
1256 => "11110111111111101111110111111001",
1257 => "11111111111101110000100111111101",
1258 => "11110100111111000000011011111111",
1259 => "00000000111111011111101000001000",
1260 => "00000001111100000000000000000101",
1261 => "00000011000000001111111000000100",
1262 => "11111011111101101111011100000000",
1263 => "11110111111100111111111011111110",
1264 => "11111111111110000000001011101011",
1265 => "11110011111011000000000011110011",
1266 => "11010001111001111111110011011110",
1267 => "11111010111101011111011011111100",
1268 => "11111011111110100000000111111010",
1269 => "00000001110110111111101111110101",
1270 => "11110110111111101110001000000001",
1271 => "11110001111100111111101111110100",
1272 => "11111111110110000000100011101000",
1273 => "11110001111010101111011011110110",
1274 => "11010101111001101111011011100110",
1275 => "11111111111010101111001111111001",
1276 => "11110001111011100000011111101111",
1277 => "00000111111011011110100111110111",
1278 => "11101111111011011110101000000011",
1279 => "11101011111101111111101111110010",
1280 => "11111010110101110000001111100011",
1281 => "11101001111011111111000011110001",
1282 => "10111001111011111111000111001100",
1283 => "11111011111100111111101111101111",
1284 => "11111111111010110000011011101100",
1285 => "00000111110011101111010111101100",
1286 => "11110100111100011110001100000000",
1287 => "11110110000000001111111011100111",
1288 => "11110101110101111111011111101101",
1289 => "11101100111010101111001111110001",
1290 => "11001000111010001111110011101010",
1291 => "00001000111101011111011011111110",
1292 => "11111010111000000000101011110011",
1293 => "00000101110001011111010111111000",
1294 => "11110000111101111101110000000101",
1295 => "11101110111011011111010011101110",
1296 => "00000001110010100000010111100000",
1297 => "11110010110111110000000011101011",
1298 => "11000101110100010000100111001110",
1299 => "00000100110111011111100100000000",
1300 => "11111010111100011111110011101101",
1301 => "11100111110011111111011011111111",
1302 => "11101110111101011110011100000011",
1303 => "11101111111011011111101111110010",
1304 => "00000001110010100000100111101110",
1305 => "11101100110110111111100111101000",
1306 => "11000110110111000000000011001111",
1307 => "11110100110110001111011011110011",
1308 => "11110011111011010000010011110011",
1309 => "11011100110111111111001111111101",
1310 => "11100100111100111110011000000101",
1311 => "11101101111111010000010111101101",
1312 => "00000100110101010001001111111001",
1313 => "11101100111000111111001111110011",
1314 => "11001111111010101111101011011100",
1315 => "11111110111000111111100111111001",
1316 => "11111100111001110000100011111100",
1317 => "11011110111001001111110011110101",
1318 => "11110101000000011111010000000011",
1319 => "11110001000011011111100011101111",
1320 => "11101101111010101111001011110001",
1321 => "11011110111001011110101111110000",
1322 => "11011000111011001101111111011110",
1323 => "11111111110111101110100111100011",
1324 => "11101101111011000000000111110110",
1325 => "11101000111001001110101011100100",
1326 => "11100011111010101111100100000000",
1327 => "11101111111100011111010011011100",
1328 => "11110101110101101111000111111001",
1329 => "11011011111001011101110111110010",
1330 => "11101111111011011101101011111110",
1331 => "00000000111010111111010111111100",
1332 => "11101100110101010000010011110010",
1333 => "11100011111100111110010111100101",
1334 => "11101011111010101111101000000001",
1335 => "11110011111100011111010111100011",
1336 => "11110111111010101111100111111010",
1337 => "11101110111110011111101111111101",
1338 => "11111000111111011111000011111110",
1339 => "00000010111100111111011011111011",
1340 => "11111010111010000000011011111111",
1341 => "11110100111101101111000011110101",
1342 => "11110011111101100000000000000100",
1343 => "11111010111110101111010111110000",
1344 => "11111111111101011111101111111101",
1345 => "11111000000000000000001000000010",
1346 => "11111101000000001111010011111100",
1347 => "00000100111111100000001111111110",
1348 => "00000010111101000000010100000011",
1349 => "00000101111111111111101111111000",
1350 => "11111010111111010000011111111110",
1351 => "11111110000000100000000011111000",
1352 => "00000000000000000000000000000000",
1353 => "00000000000000000000000000000000",
1354 => "00000000000000000000000000000000",
1355 => "00000011000000100000000000000101",
1356 => "00001011000001010000100100000011",
1357 => "11111100000001000000100000001010",
1358 => "00010001000001100000000000000101",
1359 => "00000110000001010000101100001000",
1360 => "00001111000000100000001100000001",
1361 => "00000011000001000001101100001111",
1362 => "00000001000001110000100000000010",
1363 => "00000100000001100000001000000100",
1364 => "00000100000001100000100000000101",
1365 => "11101011000000010000101000000011",
1366 => "00010011111111110000000100000000",
1367 => "00000111000000110000010000000101",
1368 => "00001000000001000000000000000110",
1369 => "00000111111111110001010100010011",
1370 => "00000110000001000000010000000010",
1371 => "11111101111101111111101011111001",
1372 => "00001010111111110000010011111100",
1373 => "11101011111111110000011100000000",
1374 => "00010001111110110000001000000001",
1375 => "00000001111110100000000100000111",
1376 => "00000000111111101111001100000010",
1377 => "00000110111111110000110000001101",
1378 => "11111011111111100000000100000001",
1379 => "11110110111111001110100111100101",
1380 => "00000001111100000000101011101111",
1381 => "11100010111011000000000111110000",
1382 => "00001111111101011111100000000011",
1383 => "11111000000000001111100111111011",
1384 => "11101011111010011110010111111001",
1385 => "11110101111010111111000000010010",
1386 => "11101101111011011111011111111111",
1387 => "11110011111101111111001111101010",
1388 => "00010110111010100000011011110111",
1389 => "11110001111011100000011111110011",
1390 => "00010001111011001111011000000101",
1391 => "11101100111100111111101111111100",
1392 => "11110001111101111111111000001010",
1393 => "11110100111101001111000100010011",
1394 => "11110011111101011111110000001101",
1395 => "00001110111011111111001100000110",
1396 => "00010110000101010000101111111000",
1397 => "00000110111111000000000100010000",
1398 => "00001110000100000000000100000011",
1399 => "11110110000001101111000000000110",
1400 => "11101010000100011111110000001000",
1401 => "11101111000010011111011000001100",
1402 => "11111100000010101111011100000110",
1403 => "00000101000011111111000011111110",
1404 => "11111111000110100000010011111101",
1405 => "11110010000010000000100100001011",
1406 => "00001111111111111111111111111100",
1407 => "00001011000111001111101111110110",
1408 => "11111110000001110001001000000000",
1409 => "00000000111111111111111000010001",
1410 => "00001000000000011111111011111011",
1411 => "00000001000010001110111000000010",
1412 => "11110010111011111111111100000011",
1413 => "00000001000000111110111100001001",
1414 => "00000101111011011111111111111101",
1415 => "00000001000011101111010100000001",
1416 => "11111000000000001111010111101010",
1417 => "00000010000000111110111000010010",
1418 => "00000100000000010000001011101011",
1419 => "11111001000100101110001011111101",
1420 => "00000011111101100000011000000011",
1421 => "00001001000000000000010000001010",
1422 => "00001110111100111111110100000010",
1423 => "11111111000110000000001000000010",
1424 => "11111111000000101111101111111011",
1425 => "11111110111111101111011100001011",
1426 => "11111101111110001111001000000001",
1427 => "11111110000001011111000111111010",
1428 => "00000011000000010000101100000000",
1429 => "11111100000001110000010000010001",
1430 => "00001101000000111111011100000101",
1431 => "00001011000010101111110000001101",
1432 => "11111010111101110000000100000100",
1433 => "11111101111111011111110100001100",
1434 => "11111111111110101110101011111101",
1435 => "11111011111111101111010011110101",
1436 => "00000111111110100000100011110110",
1437 => "11101101111101010000101000000000",
1438 => "00001100000000011111011100000001",
1439 => "11111011000000011111110011110101",
1440 => "11111110111101101111100011111100",
1441 => "11110100111101111111010000010000",
1442 => "11111010111110001111001100000100",
1443 => "11111110111100111111011011110111",
1444 => "00000111111111110000100111111100",
1445 => "11101011111110010000100011111111",
1446 => "00001011111110111111111100000010",
1447 => "11111000111101011111011000000010",
1448 => "11101101111111001111001100000100",
1449 => "11111001111111001110110100001111",
1450 => "11110111111110101111101100000010",
1451 => "00000011111110011111111011111100",
1452 => "00001011000000010000100111111100",
1453 => "11110111000000100000011100000110",
1454 => "00010000000000010000001100001000",
1455 => "11111100111101110000011000001000",
1456 => "11110110111110110000000100000101",
1457 => "11111100111110101111101000001111",
1458 => "11111101111110111111111000000001",
1459 => "00000010000000001111111100001001",
1460 => "00010111000000110000101100000101",
1461 => "00001000000100010001010000001011",
1462 => "00001110000000110000011000000110",
1463 => "00001011000001110000100000010000",
1464 => "00010110000101000000001000001111",
1465 => "00001100000001010001101000010000",
1466 => "00000101000001100000100100001111",
1467 => "00001101000010100000101000001110",
1468 => "00010000000100110000011100000110",
1469 => "00010000000011010000010000010101",
1470 => "00001100000101000000101100000101",
1471 => "11111001000100000001011000010101",
1472 => "00010111000011010000101100001011",
1473 => "00000001000011000001110000001100",
1474 => "00001110000010100000010011110001",
1475 => "11110100000100100000011100000101",
1476 => "00000000000001000000100011111011",
1477 => "11101110000001111111110000000000",
1478 => "00001110000000010000000100000111",
1479 => "00010010111101000000101000000101",
1480 => "00010001111101010000011011110011",
1481 => "00001000111111100000111000010000",
1482 => "00000101111111110000100011110110",
1483 => "11110110000110101110111111111001",
1484 => "11101010000101000000011011110110",
1485 => "11111000111111111110110111111100",
1486 => "00001110111111101111001000001000",
1487 => "00000000000011011111110111110111",
1488 => "00000000000001011111111000000101",
1489 => "00000101111110011111010000001011",
1490 => "11111000111110101111101111101000",
1491 => "11111100000111111111010100000000",
1492 => "11101011000101010000101111110011",
1493 => "00000101000011001111110100000000",
1494 => "00011010000001111111011100001000",
1495 => "00001100000001110000000111111000",
1496 => "00001001111111110000110100000010",
1497 => "00001100000000001111010100010001",
1498 => "11111001111111001111101011110011",
1499 => "00000011000110001111111011111010",
1500 => "11011000000000001111111011111110",
1501 => "00010000000000011110111100010010",
1502 => "00010000000000001111101111111100",
1503 => "11110111001110101111101111110111",
1504 => "00000010000010100000011011110101",
1505 => "11111100000000011111110100010110",
1506 => "11111000000001001111100111101010",
1507 => "11111001000111011111111000000011",
1508 => "11010010000001111110001111111111",
1509 => "00010010000000001100101100011000",
1510 => "00001110111111000000010011010010",
1511 => "00001010001010011111110000000111",
1512 => "11111010000001000001000011011000",
1513 => "00010010000000101111100000011011",
1514 => "11111110000010110000011111010101",
1515 => "11110001000101101111011111111111",
1516 => "11100101111111001110111000000001",
1517 => "00010100000000011101101100010111",
1518 => "00001100111101111111101011101110",
1519 => "11111110001010110000000100010110",
1520 => "00000010000000100000000011101010",
1521 => "00000100000000110000100000011100",
1522 => "11111011000001000000110011100000",
1523 => "11101100000011001110111000000111",
1524 => "11011100111110000000001000000100",
1525 => "00011101111110101101111000011010",
1526 => "00000100111101011111101000000100",
1527 => "11111111000101111111100100001101",
1528 => "11110111000011001111111011110001",
1529 => "00001101000000101111110100001110",
1530 => "11110100000010000000011111100111",
1531 => "11110101000001010000001000000010",
1532 => "11101110111100110000010000001101",
1533 => "00011101111101111101010100011111",
1534 => "00001001111101001111110000000010",
1535 => "00010011000100001111111000011001",
1536 => "11111010000000110000101111101011",
1537 => "00000110111111001111111100010011",
1538 => "11110110000001000000001011101111",
1539 => "11111010000001100000011000001010",
1540 => "11101101111111100000000000000000",
1541 => "00001101111111101110111100001110",
1542 => "00001100000000111111110100000001",
1543 => "00000010111111110000010100001111",
1544 => "00000111000001100000100111101100",
1545 => "00000011000001010000010100001110",
1546 => "11111100000011010000101111101001",
1547 => "11111001111110110000001000000100",
1548 => "11110001111101001111110011111100",
1549 => "11101001000000111111011111111010",
1550 => "00001100111111111111111000000100",
1551 => "11111100111111010000000100000111",
1552 => "11111110111110011111110011111111",
1553 => "00000110111111100000001000001111",
1554 => "11111100000000000000101111110011",
1555 => "11110101111101111111100011110001",
1556 => "11110101111110010000001111111111",
1557 => "11110100111010110000011000000100",
1558 => "00001001111010101111010100000010",
1559 => "11111000111101001111101100000010",
1560 => "11110001000000011111110000000010",
1561 => "11111001111111101111011100010001",
1562 => "11111010111110101111110011111111",
1563 => "00000110111110111111110111111100",
1564 => "00010100111110110000100100000001",
1565 => "11101110111110110001111000000000",
1566 => "00001101111110110000000000000011",
1567 => "11110110000011001111111100000111",
1568 => "11110100111111001111100100001000",
1569 => "11111010111110001111110100001111",
1570 => "11110111111111001111111100010001",
1571 => "11110101000001001111011011111010",
1572 => "00011010111101100000100111111111",
1573 => "11111010111111010001011000001000",
1574 => "00001100111111001111111000010110",
1575 => "11111110000001010000011100001100",
1576 => "00001001111101111111011000010011",
1577 => "11110110111110110000100000010001",
1578 => "11111100111111000000000000010011",
1579 => "00001101000010110000000111101110",
1580 => "00000100000001111111111011110101",
1581 => "11101010111110100000100011110000",
1582 => "00010000000000100000100000000111",
1583 => "00000000000001000000001011101111",
1584 => "00000000111011111111101100000100",
1585 => "00000111111101101111011100010011",
1586 => "11111101111100100000000000000011",
1587 => "00000011000100111111101111101000",
1588 => "11111100111110011111101111110110",
1589 => "11100110111100110000010011101010",
1590 => "00100001111111011111011000010011",
1591 => "11110101000001011111110111100110",
1592 => "00001111111100111111110100001001",
1593 => "11101100111011111110011100010101",
1594 => "11110010111010111110100100001100",
1595 => "00001100000011011111100011111000",
1596 => "11101000000110001111011011111101",
1597 => "00000011111111101110111100000011",
1598 => "00001100000001011111100100001111",
1599 => "00000000111011001111000111011010",
1600 => "00000101000001000001001000010100",
1601 => "11110110000000011110110000010111",
1602 => "11111110000000001111011111110100",
1603 => "11110101001001111111101011110110",
1604 => "11011001111101101110001100000101",
1605 => "00001000111100001101011000001011",
1606 => "00010001111100010000010011101111",
1607 => "11111101111111111110111111110011",
1608 => "00000011000000110000010011101101",
1609 => "00000001111111101111001000010011",
1610 => "11111000111110110000010111100100",
1611 => "11110011000110000000000111111001",
1612 => "11011110111101111110011100000110",
1613 => "00001100111110101101100000001111",
1614 => "00000010111111011111110011101011",
1615 => "00000001000110101101111011110111",
1616 => "11100101000011001111110011100110",
1617 => "00000111111110111110111100011010",
1618 => "11111110000001110000000111101001",
1619 => "11111011000110010000001111111101",
1620 => "11011011111100111110010111111110",
1621 => "00010001111101001100100000011000",
1622 => "00010010111110010000010111111100",
1623 => "11111010001001111110010111110100",
1624 => "11110001000000011111101011100001",
1625 => "00000010111111101110100100010011",
1626 => "11111011000000000000001111100110",
1627 => "11110100000001100000000100000000",
1628 => "11101011111100101111000011111100",
1629 => "00011111111111001100101000101010",
1630 => "00010110111010101111101111111101",
1631 => "00000111000010101110100100001010",
1632 => "11101111000010111111101111001110",
1633 => "00000000111111111111000000011101",
1634 => "11111111000001100000011111100000",
1635 => "00000111000001110000010100000100",
1636 => "11111111111000110000101000000101",
1637 => "00100111000000001101100100100101",
1638 => "00001100111101011111110111110110",
1639 => "11111111000100001111000000010110",
1640 => "11110111000011011110111011100010",
1641 => "00000110111110111111101000010001",
1642 => "11111100000001100000010111101011",
1643 => "11111110000001000000000011111101",
1644 => "11101100111010001111110000000000",
1645 => "00011000111111001101000000011010",
1646 => "00001010111011110000001011110011",
1647 => "00000100000000011111100100001110",
1648 => "11111101000001101110111111010100",
1649 => "00001010111100101111100100010001",
1650 => "11111011000000000000100111100101",
1651 => "00000000111111101111101111110100",
1652 => "11101011111101111111010111111000",
1653 => "11101011111100101110011000000101",
1654 => "00001111111110101111100100000101",
1655 => "00001011000000111111011011111001",
1656 => "11110110111110111110111011100011",
1657 => "11111101111111001111010000001111",
1658 => "11111001111101111111100111100100",
1659 => "11110101111010111111010111110001",
1660 => "11110001111100001111101111110111",
1661 => "11101111111111101111010100000001",
1662 => "00001011111101011111100100000100",
1663 => "11110110111011001111101000001011",
1664 => "11101011111101111111000111111100",
1665 => "11101010111101001110101000001111",
1666 => "11110100111101011111011011110110",
1667 => "11111110111111001111100011101111",
1668 => "11111100111100100000001111110010",
1669 => "11100101111100111111111111110110",
1670 => "00010010111110001111011000000100",
1671 => "11110100111111110000010000000101",
1672 => "11111000111010111110101111110100",
1673 => "11110011111100010000101000010011",
1674 => "11110111111101011111111111101110",
1675 => "11111011111111010000001011110010",
1676 => "11110110111101010000000011110111",
1677 => "11101101111101101111101011111101",
1678 => "00001000111101001111111100000110",
1679 => "00000010111111110000111100000100",
1680 => "11111101111010011111100011110111",
1681 => "11110110111101001111100100010010",
1682 => "11110110111011101111011011101001",
1683 => "11111111000011000000001011110100",
1684 => "11100101111110001110011111110100",
1685 => "11110111111100101110101011110111",
1686 => "00010001111101101111011111111101",
1687 => "11111101111111110000110000000111",
1688 => "00000110111111011111111111111000",
1689 => "00000010000000011111110100010011",
1690 => "11110001111111000000000111101111",
1691 => "11111000111111011111011011111011",
1692 => "11100000000000001110110011110001",
1693 => "11101001111100101110110011101000",
1694 => "00001111111100011111100011110100",
1695 => "11110000110110110000111011111111",
1696 => "00010101111010101111100111101000",
1697 => "11101001000001001111111000010000",
1698 => "11111101111111111111100011100110",
1699 => "00000100111011010000110011111110",
1700 => "11100111111110001111000000001000",
1701 => "11110100111111001111100011110111",
1702 => "00010000111110101111100100001110",
1703 => "11111001111000110000110011011101",
1704 => "00001110111110100000111100000011",
1705 => "11111000111111110000000100010101",
1706 => "11111000111110111111100011110110",
1707 => "00000110000001000000010111110100",
1708 => "11100100111111111110111100000000",
1709 => "11111110111101111110010011111101",
1710 => "00001111111111001111100111110111",
1711 => "11111000111111111110101011100011",
1712 => "11110010000000000000010111111110",
1713 => "11110110000000011110000000011111",
1714 => "11111101111111111111010011101000",
1715 => "11110010111101111111111000000011",
1716 => "11100110111100101110011100000010",
1717 => "11111110111111011110000100000001",
1718 => "00010111111110000000011011101001",
1719 => "11110010111110111110001111100111",
1720 => "11101101111111111111111011100110",
1721 => "11110010111110111101110100110101",
1722 => "00000001000000001111011111110010",
1723 => "11110100000000111111111000000010",
1724 => "11100100111101101101101100000011",
1725 => "00001001111111111100100100000101",
1726 => "00000010111100100000010111100110",
1727 => "11111000000010011100110011110110",
1728 => "11101111000000011111101111010101",
1729 => "11111101111111111110000101001100",
1730 => "00000110111110011111101011101100",
1731 => "11110100111110001111100100000101",
1732 => "11100110111100011111001100000110",
1733 => "00001100000010001011111100001100",
1734 => "00010011111100010000000111100001",
1735 => "00000011111101101101111011111111",
1736 => "11011111000000011111001010111110",
1737 => "00000010000000001110110100110101",
1738 => "11111111111111010000001011011011",
1739 => "11111101000000001111110000000101",
1740 => "00000100111101110000110011111110",
1741 => "00001111000000101101001100001010",
1742 => "00001110111101001111010011100000",
1743 => "11110100000001101110110100001100",
1744 => "11100111000001101110011111010100",
1745 => "11111110111101111111111000010000",
1746 => "11111111111101010000000111100001",
1747 => "11111001111111001111111011111111",
1748 => "00000100000001000000010100000100",
1749 => "00000001000011011110110000010101",
1750 => "00010011000010011111011111100010",
1751 => "00000001111111101111110000001110",
1752 => "11100100000001101111010011101000",
1753 => "11111110111110101111101100001100",
1754 => "00000100111111110000000111110100",
1755 => "11110100000000011111100111110000",
1756 => "11100110111100001110111011111000",
1757 => "11010001111101001101100011101111",
1758 => "00001110111010011111110011101011",
1759 => "11111100000000111111100111101101",
1760 => "11110100111011011110101111011101",
1761 => "00001010111011101110101100010010",
1762 => "11111001111011100000000011100000",
1763 => "11101110111010101111010011110000",
1764 => "11010000111001111110011111101011",
1765 => "11101110111000111101011000000001",
1766 => "00001000110101111111001000000011",
1767 => "11101101111000101111010011110101",
1768 => "11100010111100111110011111011111",
1769 => "11100011111010011110011000010000",
1770 => "11110010111100011110110111100000",
1771 => "11110011000000001111111011101111",
1772 => "11110110111110010000100011110100",
1773 => "11011110111111001111011011110110",
1774 => "00001111111110001111110000000010",
1775 => "11111010000000010000011100001011",
1776 => "00001111111001101110101111110110",
1777 => "11111010111100100000111100010000",
1778 => "11111100111100111111111111101111",
1779 => "11110001111101101111101111101000",
1780 => "11100111111000011111011011110111",
1781 => "11101101111101011110100011110101",
1782 => "00001001111011101111000011111001",
1783 => "00000010111100011111001111111101",
1784 => "11101011111000101111100111100011",
1785 => "00000100111001101101111100010001",
1786 => "11110011111100101111111111100000",
1787 => "11110100000010111111001011111011",
1788 => "11111101111110110000010111111011",
1789 => "00000100111110101111110000000001",
1790 => "00010010111100111110111100001001",
1791 => "11111000111111011111110111111101",
1792 => "00000010000001001111100000000001",
1793 => "11111010111101001110111100010000",
1794 => "11111011111111001110111100000011",
1795 => "11111010111000101111100111101100",
1796 => "00001000000000010000100011111101",
1797 => "11100101000000111111111111101001",
1798 => "00001011111111001111101000000111",
1799 => "11111001111000001111101111101001",
1800 => "11111100111100011111011011111100",
1801 => "11111100111010111111010100010011",
1802 => "00000001111010111111111000000110",
1803 => "00000100110011001111110011110111",
1804 => "00000100111111100000011111111100",
1805 => "11101111111110110000010011101101",
1806 => "00001110000010111111101000000101",
1807 => "11101011111011000000010111111101",
1808 => "11110111111101110000011011111011",
1809 => "11100110000001011111110100011001",
1810 => "11111101111111111111001100000100",
1811 => "11111010110010111111011011111010",
1812 => "11100111111101101111101100000100",
1813 => "11110001111111111111000111111000",
1814 => "00001101111111101111110011101011",
1815 => "11110100111001111110110111101000",
1816 => "11001011111111011111011111110011",
1817 => "11011111111111001111001000101011",
1818 => "00000000111110011111111011101011",
1819 => "11111011111011101111111100001000",
1820 => "11110010111011111110111000000101",
1821 => "00000101000000011111000000000000",
1822 => "00101011111110110000100011011100",
1823 => "11110010111011101101100111100011",
1824 => "11011010000010011111001111110001",
1825 => "11101011111111111110101001001010",
1826 => "00001000000001001111010011101011",
1827 => "11111110111111100000100000000101",
1828 => "11111001111101011101110000000101",
1829 => "00001110000000001110001000000100",
1830 => "00101000111110010000000111111101",
1831 => "00000000111100111110110011100010",
1832 => "11111000000011000000101011100000",
1833 => "11110101000001001110110001010111",
1834 => "00000101000001000000000100000001",
1835 => "00000100000000110000001111111010",
1836 => "11110010111111101101111111111100",
1837 => "11111010000000001011110011110000",
1838 => "00011100111111110000101000000010",
1839 => "00000100111101101101100011100010",
1840 => "11101011111101111111010011001011",
1841 => "00000101111111111101101000100111",
1842 => "00000110111111100000011011011111",
1843 => "11111101000001100000000011111101",
1844 => "11101111000001011111010000000100",
1845 => "11110111111110001101100111111001",
1846 => "00001111111110010000000011011001",
1847 => "00000100000001101111110100000100",
1848 => "11101111000000011111110011011100",
1849 => "11111000000000101111100000011001",
1850 => "00000000111110110000001011100000",
1851 => "00000001000000100000001011111100",
1852 => "11110111111110001111111011111110",
1853 => "00000111111011101111101100010100",
1854 => "00001101111110110000001011101100",
1855 => "11111110000000110000011100001010",
1856 => "11100100000001001111110011111011",
1857 => "00000101000010100000100000010001",
1858 => "11111111000001000000011011111011",
1859 => "11111011000010111111011111110011",
1860 => "11110101111111010000000111110010",
1861 => "11110101111000111111001111111110",
1862 => "00010000111101101111101111111001",
1863 => "11111001111111110000000000000011",
1864 => "11111101111100011111010011110000",
1865 => "00000101111101111111100100010001",
1866 => "11111100111101011111100111110100",
1867 => "11101001111100101110111111110111",
1868 => "11101111111100111111110011110001",
1869 => "11111111111001011110010100001110",
1870 => "00010000111110011110111111111111",
1871 => "11110100111100001111110000001000",
1872 => "11110110111110101101111111101100",
1873 => "11101111111001011111010100010010",
1874 => "11101110111100101111000111100010",
1875 => "11111001000001101111100111101011",
1876 => "11110101111100010000010011110011",
1877 => "11100101111110011111100011110101",
1878 => "00010001111100011111101111111111",
1879 => "11110111000000000000011000000111",
1880 => "00001010110110101110001011110100",
1881 => "11111010111011100000110000001111",
1882 => "11110111111010101111001111101101",
1883 => "11101110111101011111101011110110",
1884 => "11110010111001000000110011110101",
1885 => "11111000000000001110111000000011",
1886 => "00001011111100001111001011111011",
1887 => "00000011111100110000010000001011",
1888 => "11111000111110110000001111110101",
1889 => "00000100111100101111100000010000",
1890 => "11110101111110110000010011101110",
1891 => "11101100000010011111010000000100",
1892 => "11110100111011100000010111110111",
1893 => "11110010111110001111101011111010",
1894 => "00010011111010001111010011111110",
1895 => "11110001111111000000100000001100",
1896 => "00001111111101111110100011110000",
1897 => "11101011111101100000100000010100",
1898 => "11110001111110001111110011101101",
1899 => "11111100110110101111100111111011",
1900 => "11111101111101100000100011110101",
1901 => "11110011111100101111100111101100",
1902 => "00001101111011001111010111111001",
1903 => "11111001111110010000110100001010",
1904 => "11110010111101011111001111110101",
1905 => "11111100111110011111011000010101",
1906 => "11111000000000011111010011110011",
1907 => "11110101110010001111110100000011",
1908 => "11111110111100000000110011111101",
1909 => "11111010111110001111111011111011",
1910 => "00010001111100111111000011111111",
1911 => "11110111111101110000010000001000",
1912 => "11010100111101101110111011111001",
1913 => "11100101111101100000101000011111",
1914 => "11111000000000111111110011111011",
1915 => "11111110110100111111011100000011",
1916 => "11110001111111100000001000000100",
1917 => "11111100000001101111011111111001",
1918 => "00000100000000011111110111100110",
1919 => "11111000111110011111000100000001",
1920 => "10011010111110101111100111111110",
1921 => "11100111000000001111001000110110",
1922 => "11111001000001011111101111100000",
1923 => "00000000111101100000001000010001",
1924 => "11011111111110111110011000001010",
1925 => "00010001000010101101111000001100",
1926 => "00100111000000000000011011010010",
1927 => "00001011111111011110110100000110",
1928 => "11010101000001011111111011011111",
1929 => "00000001000000101111010100100101",
1930 => "11111101111111110000011111100011",
1931 => "00000101000001111111110000001000",
1932 => "11101000111110101101010000000111",
1933 => "00010010111111011011111111110111",
1934 => "00101011000000000000011011110011",
1935 => "11111100000000101110000111011000",
1936 => "00000011000010101111110011011111",
1937 => "11111110111110001101110000111000",
1938 => "00001000111111001111111111011100",
1939 => "00000001000010001111101111110110",
1940 => "11111010111101001111010100000000",
1941 => "00000101111101001101100011111110",
1942 => "00001111111011111111111000001110",
1943 => "00001001000001111100111111110110",
1944 => "11111001000001001111001111101100",
1945 => "00000011111101101100110000011000",
1946 => "11111110000000100000100011101101",
1947 => "00000001000001000000001000000101",
1948 => "00000011000001000000010011111100",
1949 => "00010111111100010000001000011001",
1950 => "00000111000000111111101000011010",
1951 => "11111111000001111101110111111101",
1952 => "11110000000010010000011000001001",
1953 => "00000010111111101101111000010100",
1954 => "11111011000010001111111011111111",
1955 => "11111111000000111111010111111011",
1956 => "00000110000000010000011100000000",
1957 => "11101011111101011111111100001001",
1958 => "00000110000000111111111111111001",
1959 => "11111101000010111111001111110110",
1960 => "11111000111111000000001000000100",
1961 => "00000101111111111110010000010010",
1962 => "11111101111110011111110000000000",
1963 => "11110101000000101110110011101100",
1964 => "11111101111111100000110111110010",
1965 => "11111010111101000000001100001011",
1966 => "00001111111110111111101000000000",
1967 => "11101110111111100000001000001000",
1968 => "11110101111111101111101100000001",
1969 => "11111101111011111110100100001110",
1970 => "11111000111011111111010111111110",
1971 => "11110101111010001111000111100101",
1972 => "11101000111010101111100111110011",
1973 => "11111011111101011111001000001001",
1974 => "00001101111100101111000100001001",
1975 => "11111001111001101111101100000010",
1976 => "11100111111110111111001111110101",
1977 => "11110001111001001110000100001110",
1978 => "11110001111100001110111111101010",
1979 => "11101011111111101111100000000001",
1980 => "11110101111110100000010111110100",
1981 => "11111111111110101101111000000100",
1982 => "00001100111101001111100100000010",
1983 => "11111011111111110000101000010000",
1984 => "00001001000001001110010111111110",
1985 => "11111001111110110001100000010011",
1986 => "11110111000000101111110111111100",
1987 => "11101110000110011111101111111000",
1988 => "00000111110111000001010111111011",
1989 => "00000001111110010000000100001100",
1990 => "00001110111100101111011000001101",
1991 => "00000110000101100000001000001101",
1992 => "00001100000010001111111000000001",
1993 => "00001010111011110001101000001110",
1994 => "11101110111110001111101100000010",
1995 => "11101111000010011110011011101011",
1996 => "11111110110101100000111100000010",
1997 => "11101001111101001111100111101001",
1998 => "00001010111101001110111111110100",
1999 => "11100110000010011111000111110110",
2000 => "11110101111011111101001011101100",
2001 => "11111010111001001110101100001111",
2002 => "11101110111011000000000111110110",
2003 => "11110100111010111111111000000100",
2004 => "00000110111011110000001111111100",
2005 => "11111111000001111111110100000000",
2006 => "00000110111110011111010111111011",
2007 => "11110110111110001111110100010100",
2008 => "11110100000001001111110111111100",
2009 => "11111100000010000000010000010101",
2010 => "11110101000000011111111000000001",
2011 => "11110001111101001111001011111001",
2012 => "00000010111000110001101111110111",
2013 => "11110010111111101111011111110100",
2014 => "00001010111100001110111111111011",
2015 => "11101010000010110000001000001100",
2016 => "11010110111100001110010111110100",
2017 => "11110001111100000000000000011110",
2018 => "11101011111101111111101011110011",
2019 => "00001000111010100000001100001100",
2020 => "11100010111101001111110100000110",
2021 => "00010011000000001110101100010101",
2022 => "11111111111111010000010011100101",
2023 => "11111110000011001110010000011001",
2024 => "10000001000010100000110011111011",
2025 => "11101011000011101111100000011001",
2026 => "11110101000100100000001111010111",
2027 => "11111011000000010000001000000111",
2028 => "11011001111010011111000000001000",
2029 => "00100001000001011101101100010111",
2030 => "00010101111101010000011111110001",
2031 => "00000110000010001100011111111011",
2032 => "11011101000100011111110111101010",
2033 => "00001011000001111110110100011101",
2034 => "00000011000010110000010111101010",
2035 => "11111111000101000000010011111110",
2036 => "11110001111100001110110100000001",
2037 => "00011011111110101101100000010010",
2038 => "00100011111011110000000100010000",
2039 => "00000111000010101101010011010100",
2040 => "00000000000101101111101011101011",
2041 => "00000111111110101100100100011001",
2042 => "00000101000000010000000111111001",
2043 => "11110100000011101111011111111110",
2044 => "11110010111011001111011111111001",
2045 => "00001101111100001101001100010110",
2046 => "11111110111011001111000000010001",
2047 => "00000010000011101101010111110001",
2048 => "11101110000010001111011111100111",
2049 => "00000100111011111100111000000111",
2050 => "11110101111111010000010111101101",
2051 => "11111010111101011111111011110101",
2052 => "11110110111100011111111111111100",
2053 => "00010001111110011111010000011001",
2054 => "00001101111111101111000000011111",
2055 => "11111100111110011110101111111011",
2056 => "11100010000010011111111111111100",
2057 => "11111010111100001110101000010001",
2058 => "11110100111111000000000011111000",
2059 => "11111100111101011111110111101011",
2060 => "11110101111101111111011111111000",
2061 => "11101010111101111111100000000010",
2062 => "00001100111101001111011100000110",
2063 => "11111000111111101111001000001010",
2064 => "11101101111101010000011011111111",
2065 => "11110101111101111101011000001111",
2066 => "11110100111101101111011111111111",
2067 => "11110100111001111111111011110111",
2068 => "11111101000000101111111111110100",
2069 => "00000100111100111111001011111111",
2070 => "00001101111101011111000000000001",
2071 => "11100101111011001111100100000101",
2072 => "11101100111100111111100111111011",
2073 => "11101011111111111110011100010011",
2074 => "11111010111110011111010011111011",
2075 => "11100100111111101110110011110010",
2076 => "11101011111101100000001011110011",
2077 => "00001011000001001110110000001010",
2078 => "00010001111100101111000000000011",
2079 => "11101000111100100000111000001010",
2080 => "00000011111111011110001111110100",
2081 => "11101110111011000000111100001101",
2082 => "11110111111110001110111011100110",
2083 => "11110100000010000000001011111100",
2084 => "00001100111101010000100000000011",
2085 => "11110111000001110000111100000100",
2086 => "00010000111100111111111100001000",
2087 => "00000001000011110000100000000101",
2088 => "00001010111111101110111111111011",
2089 => "00000011000000010001111000001111",
2090 => "11111100111101110000001100000101",
2091 => "11101010111111111111010111110001",
2092 => "00001111111100010001101011110001",
2093 => "11111001111101010001000111111101",
2094 => "00001110111010101111110000000111",
2095 => "11101001000111010000100000000110",
2096 => "11110110111101001101111011110101",
2097 => "11110110111100101110100100001110",
2098 => "11110010111100011111011011110010",
2099 => "11011111111101011110101011111110",
2100 => "11101101111011000001011111111010",
2101 => "11011111111100101110111011101001",
2102 => "00001110111001001110110111110111",
2103 => "11011111000011100000000100000110",
2104 => "11110000111010101110010011100011",
2105 => "11101101111110011111101100010100",
2106 => "11110110111110101111000111110000",
2107 => "11110111110100111111100011111011",
2108 => "00001101111010010001000011111110",
2109 => "11110011111110110000110011110111",
2110 => "00010011111110101111011100001010",
2111 => "11101101111000001111101011111001",
2112 => "11110001111101101110111011111110",
2113 => "11101100111101101111011100010010",
2114 => "11111001111101011110111000000111",
2115 => "11110101000010011110111111111101",
2116 => "00000010110111000001100111110101",
2117 => "11111101111101111111100011110111",
2118 => "00001100111100101110100111110000",
2119 => "11110100000111011111111000001000",
2120 => "11101011111111001110100111111000",
2121 => "11111001111100011111010100100111",
2122 => "11101111111100111111001011110010",
2123 => "11110010111000010000000011111010",
2124 => "11011101111001111110111000001011",
2125 => "00001101000000011101100100010001",
2126 => "00011000111111011111110011111101",
2127 => "00000000111111101100100111101010",
2128 => "10101100000011011111011111111001",
2129 => "11110101111100111110100000100110",
2130 => "11111101111110110000001011011111",
2131 => "11111110111111000000010000000011",
2132 => "11100010111010011111111011111110",
2133 => "00011010000010101110000000001100",
2134 => "00011001111111100000011000010110",
2135 => "00000111000011001100001011101010",
2136 => "11100100000101011111101011101101",
2137 => "00000010111111101100010100100100",
2138 => "00000010111111101111101011100110",
2139 => "00000010000101000000010111111101",
2140 => "11110111111100011111110011111111",
2141 => "00001010111100001101110011111101",
2142 => "00010000111101100000000100001100",
2143 => "00000101000110001100110011110111",
2144 => "11110110000010001110111011100100",
2145 => "00000111111101101101100100101111",
2146 => "00000000111110110000011111110111",
2147 => "11111001000001101111110111110110",
2148 => "11101000111100101111000111110000",
2149 => "00000001111000001101011000010001",
2150 => "00000101111011011111001100000010",
2151 => "11111100000010011101110000000101",
2152 => "11110000111110011111111111011001",
2153 => "11110011111101101101011100011111",
2154 => "11110010111110011111110011011010",
2155 => "11110011111011111111000111111000",
2156 => "11100111110101001111010000000000",
2157 => "11111000110111111110000100000010",
2158 => "00010011110101101110100111111010",
2159 => "11110100111011101111110111111001",
2160 => "11110011111110111110010111011111",
2161 => "11101110111011101111110000010110",
2162 => "11110100111110001111011111100000",
2163 => "11110000111011101110111011111011",
2164 => "00000000111000000000110011101110",
2165 => "11010101111001100000001111100110",
2166 => "00001101111011011110110000010100",
2167 => "11101001111100010000000011111001",
2168 => "11110111110110101110011111111101",
2169 => "11101100111010111111010000001111",
2170 => "11110111111010101110110111111010",
2171 => "11111111111100011111100111111111",
2172 => "00000010000001000000011011110101",
2173 => "00000001111110100000000100001010",
2174 => "00010001000001011111101100010000",
2175 => "11110110111001110000010100000101",
2176 => "11111011000000111111100000000110",
2177 => "11100111111110000000000100010000",
2178 => "11110100111101101110111111111011",
2179 => "11111110000001101111101111111001",
2180 => "00001000000000000000110000000000",
2181 => "00000011111110110001010100000011",
2182 => "00001101111101101111111000001000",
2183 => "11111010000010010000011111111101",
2184 => "00000011000001101111100000001010",
2185 => "11110101111111100000010000010000",
2186 => "11111101111111101111101011111111",
2187 => "11111000000001001111110011101110",
2188 => "11111011111100010000101011111010",
2189 => "11100001111111001111111011110111",
2190 => "00001110111110001111101011111011",
2191 => "11111110000100010000011100000111",
2192 => "00000111111010101111000111110101",
2193 => "11111111111100110000110100010010",
2194 => "11110011111100010000001111110011",
2195 => "11101100111011111110101011101101",
2196 => "11111111111001100000111111110011",
2197 => "11011011111001111111010011100100",
2198 => "00010011111010011110111000000111",
2199 => "11100001000000101111011011101000",
2200 => "11011111111100111101100111111001",
2201 => "11101100111010011110000100010010",
2202 => "11110001111011101111010011111100",
2203 => "11101101110011101110111111111001",
2204 => "11111011111001100001101011111001",
2205 => "11110011111110011111011011110011",
2206 => "00001110111101101111010011111011",
2207 => "11100010000000001111011000010011",
2208 => "11100010111001111111100011101001",
2209 => "11100010111110111110000100010011",
2210 => "11101011111100101110110111110100",
2211 => "11110100101111110000000100001101",
2212 => "00000000111000110001101111111100",
2213 => "11111010111101001111101111111001",
2214 => "00001001111101111110101111111110",
2215 => "11101011111101100000011100011100",
2216 => "11111010111101101111000111101111",
2217 => "11110100000001000000010100100000",
2218 => "11101101111111001111001011111111",
2219 => "11110001111001111111011000000000",
2220 => "11100101111010100000100111111110",
2221 => "11111010111110111110010011110110",
2222 => "00011010111011101111001111110011",
2223 => "11101010111111010000010111111110",
2224 => "00000100111111001110011011101111",
2225 => "11101111111101100000001000100110",
2226 => "11110101111101101111001011101000",
2227 => "11110100111000000000011100000000",
2228 => "11010011111010101110111111111111",
2229 => "00000000111111011101100011111001",
2230 => "00110000111101001111111000001011",
2231 => "11111001111101111111111011001010",
2232 => "11101110111110111111101111101011",
2233 => "11101101111101101110101001000011",
2234 => "11111110111110101111011011011010",
2235 => "11111001000001000000011000000011",
2236 => "11111101111001110000101100000000",
2237 => "00011000111110001111001000000101",
2238 => "00100110111101110000000000100100",
2239 => "00000011000000101110010111100100",
2240 => "11101100000110010000001011110101",
2241 => "00000001111101101101011100111010",
2242 => "00000000111111001111110111111110",
2243 => "11111110000010011111100111110111",
2244 => "00000010111100101111111011111011",
2245 => "11110000111011111110100111101001",
2246 => "11111010111110100000011000000100",
2247 => "00000000000100011111001000001100",
2248 => "11111110111111001110101111110011",
2249 => "00000100111101111101010100111110",
2250 => "00000100111010111111110100000010",
2251 => "11111000111101011111101011111100",
2252 => "11101000111010101101110011111100",
2253 => "00000110111110111101101100000010",
2254 => "00000111111011111111110000001101",
2255 => "00000001111101000000000011110110",
2256 => "11111110000001011111000111101101",
2257 => "00000000111101111111001100010111",
2258 => "11111001000000011111111011110111",
2259 => "11111101111110011111110011111000",
2260 => "00000000111111000000011111111110",
2261 => "11100101000001001111000011101110",
2262 => "00001101111101111111011100010100",
2263 => "11110100111111010001000100000111",
2264 => "00001100111100001111010011110111",
2265 => "11110101000000010000100000001101",
2266 => "00000001111110101111011111111011",
2267 => "00000000111111001111111000000001",
2268 => "00001001000000000001100111101101",
2269 => "11100001000000110000110011101001",
2270 => "00010011000001011111010100011100",
2271 => "11101011111101110001001000000100",
2272 => "00010000111011010000001000001000",
2273 => "11110000111111100000010000001101",
2274 => "11111111111110111111010100001011",
2275 => "00000111111110101111110100000001",
2276 => "11110111000010010000000000000010",
2277 => "00001011000001101111101000010000",
2278 => "00001100000001001111111100001101",
2279 => "11111101111010000000110100001010",
2280 => "00000010000001010000111000001000",
2281 => "11110101000011110000011000010010",
2282 => "11111011000000010000000111111010",
2283 => "11111110000010101111111100000001",
2284 => "11110010111111011111101011111110",
2285 => "00000100111101101110101100001100",
2286 => "00010011111100001111110000000010",
2287 => "00000101000000100000101100000000",
2288 => "00001000000001011111101011110010",
2289 => "11110110111111000000100000001100",
2290 => "00000001000000111111111111110011",
2291 => "00001000000000110000001111111101",
2292 => "11101111000001000000011011111011",
2293 => "11111101000000011110111000000101",
2294 => "00010000000000101111110100000001",
2295 => "11111100000001010000011000001100",
2296 => "00000110111110100000001011101011",
2297 => "11111100000000000000011100010000",
2298 => "11111010000000001111100111101000",
2299 => "11100010000001001111110000000001",
2300 => "00000011111001000000100111110000",
2301 => "11101100000000111110010111101110",
2302 => "00010001111011001110111111111100",
2303 => "11111010000001010001100000010010",
2304 => "00011100111011110000000011101000",
2305 => "11111010111110100001010100010010",
2306 => "11111011111101111111000011111011",
2307 => "11101010110011011111010100001101",
2308 => "00010000111110100001100011111001",
2309 => "00000000000010000000100111111111",
2310 => "00000100000000001111001100000110",
2311 => "11101100111001000001101100101001",
2312 => "11110110111111101111110100000001",
2313 => "11110000000000110001101000001100",
2314 => "11111000111111010000000000001100",
2315 => "11111101101101001111110100000110",
2316 => "00010101111100100001110111111101",
2317 => "11110101000010100000100011111101",
2318 => "00001000000000011111010111111110",
2319 => "11110001111010100001100100001011",
2320 => "00000010111110101110100000001000",
2321 => "11101101111100000001011100010010",
2322 => "00000100111101111111101100010011",
2323 => "11110011111000101111100100000100",
2324 => "00000110111011100000111011111011",
2325 => "11111010000010001110011011111010",
2326 => "00001110111111011111111111101001",
2327 => "00000001111100000001001111110011",
2328 => "00001010111110011110100011101111",
2329 => "11111010111011010000101000101101",
2330 => "00000011111110101111111011111000",
2331 => "11110100111011101111101000001010",
2332 => "00000011111010100000000111111011",
2333 => "00000010000010111110011000000001",
2334 => "00110000000000011111111011111011",
2335 => "11111101111100110001110111110010",
2336 => "00000110000000101110010011111000",
2337 => "11101010111001010000000001000101",
2338 => "00000110111110011111010011110111",
2339 => "11110111111011110000001100001011",
2340 => "11110001111010111111010011111110",
2341 => "00001110111111011110110100000001",
2342 => "00110001000000110000011100001110",
2343 => "11111000111110010000101011100010",
2344 => "11110111000010001110101111111001",
2345 => "11111011111011101110101101010101",
2346 => "00000111111100101111101011110111",
2347 => "00000100111110110000000011111011",
2348 => "11110000111111011101111111111011",
2349 => "11011010111101011110000111011010",
2350 => "00100101000000000000010111111101",
2351 => "11110011111011111111011011101100",
2352 => "11111100111100111111011011110001",
2353 => "11110101000001001110101000110101",
2354 => "00000011111110011111110011110011",
2355 => "00000100111101101111111011111001",
2356 => "11111110111110111110011000000001",
2357 => "11101000111111111111010111011111",
2358 => "00010110000000100000011100001010",
2359 => "11111001111001110000100011110001",
2360 => "00001111000000111111100111111111",
2361 => "11111110000001000000000100011100",
2362 => "00001000111100111111110100000011",
2363 => "00000010000011101111101000000111",
2364 => "00001001000010101111101011111011",
2365 => "11001100111111100000010011011110",
2366 => "00010100000010000000000100001001",
2367 => "00000000111111110001000111110100",
2368 => "00011100111101000000000100001100",
2369 => "11101101111100000000011100011011",
2370 => "00000010111100101111001100001000",
2371 => "00000111000000011111011000000101",
2372 => "00000100000011101111111111111010",
2373 => "11100110000000110000101111111000",
2374 => "00010011000001110000000100001001",
2375 => "11110111111110000000111111110101",
2376 => "00010011111111000000111100001111",
2377 => "11110011111110110000011100010011",
2378 => "00000100111100111111011100000110",
2379 => "11111010111100111111000100000011",
2380 => "11111110000011101111111000000010",
2381 => "00000100000010001111100100001111",
2382 => "00010000000001000000001100001001",
2383 => "11111101111011000000001111101111",
2384 => "11111100000000011111111100000001",
2385 => "00000011111101011111011100001010",
2386 => "00000110000001111111100111111110",
2387 => "00000011000011100000001011111111",
2388 => "00000100000010100000110111111101",
2389 => "00000100111110000000011000001101",
2390 => "00001001000011101111111100000101",
2391 => "00000100000001000000100011111111",
2392 => "00010011000000100000100000000100",
2393 => "00000000000001101111111000001011",
2394 => "00000110000001000000001000000100",
2395 => "11110101000001111111100111111111",
2396 => "00000011111111000000010011111110",
2397 => "11111000111110100000100011111101",
2398 => "00001100111101011111110000000000",
2399 => "00000001000001111111110000000110",
2400 => "11111100111110011111000100000001",
2401 => "11111010000001010000000000001101",
2402 => "00000010111111110000000011111110",
2403 => "00000010000000001111111000000001",
2404 => "11111011000100100001000100000100",
2405 => "11111010000001010000000100000001",
2406 => "00001011000000110000001000000101",
2407 => "00000001000001110000001100001011",
2408 => "11111110111110110000011100000011",
2409 => "00000001000000101111110000001100",
2410 => "00001100111111110000001111111101",
2411 => "11110101111111011111010100001001",
2412 => "11111111111101010001101000000100",
2413 => "11111001000000010000010111111101",
2414 => "00001011111101011111011111111111",
2415 => "11111010000110000000011000010000",
2416 => "11111101111111111110110111111110",
2417 => "00001000111111010000110100010101",
2418 => "11111010111111110000000000000101",
2419 => "11110001111111011111100100001001",
2420 => "00001001111111000001101111111110",
2421 => "00000111000000100000100100000011",
2422 => "00001111111101101111011111111100",
2423 => "11110000000010110000100100000001",
2424 => "11110111111111111110111100001000",
2425 => "11110110111011000000011100010010",
2426 => "00000000111101111111101000001000",
2427 => "11110011111111001111101000000100",
2428 => "00000010111001110001001111111010",
2429 => "00000111000001101111011000000110",
2430 => "11110101111111001111010011111010",
2431 => "00000010000011100000001011101101",
2432 => "11110110111110101110101111111101",
2433 => "00000010111001011111111000011110",
2434 => "11111101111110001111111111111101",
2435 => "11111100111110100000010011111100",
2436 => "11110001111110001111010111110101",
2437 => "00000100111111111110100011111010",
2438 => "00001101000000011111110000001001",
2439 => "11111001111111111110001111011110",
2440 => "11100110111111001111001100000011",
2441 => "11111000111011011101001100101101",
2442 => "11111101000000001111011111110010",
2443 => "00001001111101000000011111110100",
2444 => "11101101111110111110001111111100",
2445 => "11111001000001011110111011111001",
2446 => "00101100111111000000100100001101",
2447 => "11111001111011101101011111001101",
2448 => "00000000111100111111100011111101",
2449 => "11110001111111111100101000110101",
2450 => "00000011000000011111011011110001",
2451 => "00000000111111100000100011101010",
2452 => "11111011111101101110111111111000",
2453 => "11011111111110010000000111011101",
2454 => "00011100111100101111111100010011",
2455 => "11110100111101011111010110110111",
2456 => "00010001111110011111011000000010",
2457 => "11110011111101111101001000011000",
2458 => "11111110111101001111100000000100",
2459 => "00000001111111000000110011111111",
2460 => "00001100000000010000000011111001",
2461 => "00001011000001110000111000001001",
2462 => "00001110000010101111111100100100",
2463 => "00000100000000001111111111101101",
2464 => "00001110000001010000000000010110",
2465 => "00000000111111001111001000011000",
2466 => "00000001000001000000010100010000",
2467 => "00000100000010110000001100001010",
2468 => "00001000000010010000010011110100",
2469 => "11100101111101010000011011111101",
2470 => "00001101000001010000001000100010",
2471 => "11111010111110010000100011011011",
2472 => "00010101111110001111101000001101",
2473 => "11110110111100011111110000010100",
2474 => "11111100000001000000000000001100",
2475 => "00000011000001110000001011111101",
2476 => "00000111000011000000110011111011",
2477 => "11111101111111000000111111111101",
2478 => "00010011000001011111011100011011",
2479 => "11111000111111110001101111110110",
2480 => "00011011111110010000110000010011",
2481 => "00000001000000100001001100001101",
2482 => "11111010000000101111110100001100",
2483 => "00000111111010111111110111110111",
2484 => "00000101000000010000011100000001",
2485 => "00001001111100000000101100001101",
2486 => "00001100111111001111101100001100",
2487 => "11111111111101001111010000000100",
2488 => "11011111000001000000110000001110",
2489 => "11111000000010111111100100010100",
2490 => "11111000000000011111101100001001",
2491 => "00000011000001111111111000000011",
2492 => "00000100000001110001001111111111",
2493 => "00010100000010010000111000001011",
2494 => "00001110000010100000010100001000",
2495 => "00000001000000100000100000010010",
2496 => "00000100000010000000001000010000",
2497 => "00000001000001000000100000010000",
2498 => "00000101000000001111110100001000",
2499 => "11111011111111111111111011111010",
2500 => "11111001000000000000001111111101",
2501 => "11101110000000001111110011111010",
2502 => "00001110111110111111100011111111",
2503 => "11111111000001110000001100001000",
2504 => "00001010111101011111111111110010",
2505 => "00000000000000010000110100010000",
2506 => "00000010000000001111111011101101",
2507 => "11111111111111010000000011111011",
2508 => "00000011111101110000110000000010",
2509 => "00000010000000000000100000001010",
2510 => "00010101111111111111111100000100",
2511 => "00000011111111110000011111110111",
2512 => "00001000000000111111101100000110",
2513 => "00000001111101110001001000001111",
2514 => "11111011111110110000001000000101",
2515 => "00000011000100111111111100000011",
2516 => "00000101111110000000010000000101",
2517 => "11111010000000000000000011111101",
2518 => "00001000111111011111010111111111",
2519 => "11111011000111010000010100010011",
2520 => "11101100000001111111100100000000",
2521 => "00001011111110111111010100010000",
2522 => "11110111111101110000011100000010",
2523 => "11111001000101011111110000001011",
2524 => "11111000111111111111110011111101",
2525 => "00010001000001011111011000010001",
2526 => "00001100000000011111010011111101",
2527 => "11110101000001011111101000010011",
2528 => "11101111000001011111000111111000",
2529 => "11111011111110010000001000010011",
2530 => "11111011000001001111111111111010",
2531 => "11111100001001100000001111110101",
2532 => "00000100111111100000011100000011",
2533 => "00001110111110101111101000001001",
2534 => "00000101111101000000000000000011",
2535 => "00001000000011011111100011110010",
2536 => "11110001000010101111100011111010",
2537 => "00000101111101001110111000001111",
2538 => "11111100000010001111100100000001",
2539 => "11110001000100011111111111110110",
2540 => "00000001000001101111110011111011",
2541 => "00001100111110101111001100010010",
2542 => "00010010111111101111100100000100",
2543 => "00000100111110101110101011010101",
2544 => "00000110000000001111111000000000",
2545 => "11111110111110001101101000001110",
2546 => "11111100000001001111110111111111",
2547 => "11111101000011110000001111110000",
2548 => "11111010000001001111010000000001",
2549 => "11110101111101111111011100000101",
2550 => "00011001111111101111110100001010",
2551 => "11111100111100111111010111100111",
2552 => "00001010000001101111111011111101",
2553 => "11111010111100111101011000010000",
2554 => "00000011111110100000001111111011",
2555 => "11111101000011010000001111101010",
2556 => "00000011000010100000010111111010",
2557 => "11111011111100000000001000000011",
2558 => "00010110111110100000000000001001",
2559 => "00000001000000011110110000000000",
2560 => "00000101000000100000011011111110",
2561 => "11111001111111001110100100010010",
2562 => "00000110111111001111110100001001",
2563 => "11111101111111101111111000000001",
2564 => "00001000000010010000000000000010",
2565 => "00100010000011000000001000011110",
2566 => "00010011000000001111111100001011",
2567 => "00010100111100000000110011110111",
2568 => "00000010000110100000110000000011",
2569 => "00010011000000000000010100001111",
2570 => "11111101000010011111110100000110",
2571 => "11110101111111111111110000000011",
2572 => "00000100000000101111101100000001",
2573 => "11110100000001111111100000000101",
2574 => "00010000000000001111111000001100",
2575 => "00001010111110100000001000000011",
2576 => "00000010000000001111101000000011",
2577 => "00001110111101110000011100010011",
2578 => "00000100111110000000010000000110",
2579 => "00001001000011010000011111111111",
2580 => "00000001000011010000101111111001",
2581 => "11110111000000110000001000000101",
2582 => "00001111000001111111100100000011",
2583 => "00001001000001110000000100001001",
2584 => "00000110111110010000110100000000",
2585 => "00000100000100000000011000001111",
2586 => "00000001000011011111111100000010",
2587 => "11101111111010011111001011110110",
2588 => "11101101111010011111010011111001",
2589 => "11110101111101011110101111111101",
2590 => "00010010111101111110111100000010",
2591 => "11110001111010011111111111111001",
2592 => "11111000111101011110000111101110",
2593 => "11101111111001001111110000001101",
2594 => "11110101111011011111101011100111",
2595 => "11111100111101010000000000000000",
2596 => "00000011111110100000110100000111",
2597 => "00001101111110110001001000001100",
2598 => "00010000111101001111111000001001",
2599 => "11111100000000111111111100010001",
2600 => "11110110000011100000010100001010",
2601 => "11111110000001000000111000001101",
2602 => "11111101000001110000001000001001",
2603 => "11111100000000110000000100000000",
2604 => "00000000000000010000010100000010",
2605 => "11110001000001011111111000000001",
2606 => "00001011000001001111111000000001",
2607 => "00000101000000110000011000001011",
2608 => "00001110111110110000010000000010",
2609 => "00000101000001010001001000001100",
2610 => "00000101000001010000001000000000",
2611 => "11111100000000111111101111111000",
2612 => "11101000111111111111100111111011",
2613 => "11011111111110111110101011110100",
2614 => "00001111111111111111111011111010",
2615 => "11111010111101110000100100001110",
2616 => "00001010111011011111100111101111",
2617 => "11110111111111100000100100001100",
2618 => "11111111000000011111111111100001",
2619 => "11110010111110011111001011110011",
2620 => "11101101111111011111010111111010",
2621 => "11111001111101001110101100000100",
2622 => "00001110111110001111010111110111",
2623 => "11111101111110100000101000001010",
2624 => "00001001111101001111100011100011",
2625 => "11111110111111000000011000001111",
2626 => "11110110111100011111001011100101",
2627 => "11111000111101101111001111110101",
2628 => "00000000111110101111101100000110",
2629 => "00000101111110011111100100010001",
2630 => "00010100111110011111100100000000",
2631 => "11111010111101100000100000000010",
2632 => "00000111000000111111010111111101",
2633 => "11111011111100011111001100001111",
2634 => "11110111111110001111111111111000",
2635 => "11111011000010011111111111101101",
2636 => "11110101000001010000101111101010",
2637 => "11011000111101010000001011110000",
2638 => "00001111000000101111010100000000",
2639 => "11111000000000100000100100001111",
2640 => "11111110110111010000000011110010",
2641 => "11111110000000011111101100010101",
2642 => "11110011111100001111000111110100",
2643 => "00000000111010100000011111101010",
2644 => "11111010111100001111110100000100",
2645 => "11110110111010011111110000000010",
2646 => "00010011111001001111001000001001",
2647 => "11111010111110100000100000001100",
2648 => "11101101111111111111111000000001",
2649 => "11110011000000100001000000001100",
2650 => "11101110000001000000000011111010",
2651 => "11110100000000001111011011101110",
2652 => "11110111000001001111110011110001",
2653 => "11100101000011101111010111111001",
2654 => "00001100000001101111011000000100",
2655 => "11110000000001000000010100000101",
2656 => "00000010111010001111000111110111",
2657 => "11110001111111100000001100001111",
2658 => "00000010111101111111101111110100",
2659 => "11101101111111101110110111110110",
2660 => "11110010111010101111011011101011",
2661 => "11100001111011011111010111111001",
2662 => "00010010111010111111000111111100",
2663 => "11111001111111100000101000001010",
2664 => "00001001111000101110111111101101",
2665 => "11110101111010111110111100001010",
2666 => "11101101111010111111001111101010",
2667 => "11111110111000000000010011111011",
2668 => "11101110110101111111011111111011",
2669 => "11111011110110001111110000000111",
2670 => "00010110110101101111100000010000",
2671 => "00000001111001100001000100001000",
2672 => "11011110111011000000011100000010",
2673 => "00000011000000000000110000010110",
2674 => "11100111000001010000000011110101",
2675 => "11111101111100011111111011110110",
2676 => "11110110111100010000000011111001",
2677 => "11101111110111100000000111111110",
2678 => "00010011111001111111110100010100",
2679 => "11111101111110000000010000010001",
2680 => "11011101111011111111011011111111",
2681 => "00000010111101010000111000010011",
2682 => "11111001000001111111110111111100",
2683 => "11111111111111010000010111111101",
2684 => "11111011111100100000001011111000",
2685 => "11110000111001101111111011111000",
2686 => "00001011111010001111101000001010",
2687 => "11111110111111100000001100010001",
2688 => "11101110111101000000000000000010",
2689 => "11111011000001000000000100001110",
2690 => "11110100000000111111111011111011",
2691 => "11101111111101001111001000000011",
2692 => "11110000111110001111111111111100",
2693 => "11111101111101101110011011111001",
2694 => "00001011111011101111110011111111",
2695 => "11111001111010010000000000001010",
2696 => "11110111111111001110101011101101",
2697 => "11110011111001110001001000001111",
2698 => "11111001111111111111100011101011",
2699 => "11110110111101001111010011111111",
2700 => "11111010111111110000010100000100",
2701 => "11111011111111111111101100000100",
2702 => "00001011000000000000010100001000",
2703 => "11111011111101010000011000000110",
2704 => "11111100000001011111001011111011",
2705 => "11111011111101100001001000010010",
2706 => "11111110111110100000000111110101",
2707 => "00000000000000000000000000000000",
2708 => "00000000000000000000000000000000",
2709 => "00000000000000000000000000000000",
2710 => "11111111000000111111111111111101",
2711 => "11111100111111111111110011111100",
2712 => "00000110111110111111100000000100",
2713 => "00000101000000100000001011111110",
2714 => "00000000000000111111101011111110",
2715 => "00000001000000010000000111111100",
2716 => "11111110000000101110010100000011",
2717 => "00000011111111001111110111111101",
2718 => "11110100000000011111101011111010",
2719 => "11111101111110001111100111111001",
2720 => "11111110111101101111101011111100",
2721 => "00000001111110001111101000000010",
2722 => "00000000000001001111110111111111",
2723 => "00000010111110101111011011111101",
2724 => "00000010111111011110100011111110",
2725 => "11111100111111000000000011111101",
2726 => "11110111000000111111011111111101",
2727 => "11111010111110111111100111111011",
2728 => "11110111111111000000000111111011",
2729 => "00000101111101111111111011111101",
2730 => "11111001000000101111011111110100",
2731 => "11111101111110101111101000000010",
2732 => "11111001111101111111010000000110",
2733 => "11111111111111011111010100000010",
2734 => "00001001111100100000101100000110",
2735 => "11111100000100101111100000000100",
2736 => "00010001000001100000001000010001",
2737 => "11111110000011000000001000000110",
2738 => "11111001000011001111000100000011",
2739 => "11110101000110010001010000000111",
2740 => "11111100000010101110111100000001",
2741 => "00000111000010101111111000000111",
2742 => "00001001000101101111101100001111",
2743 => "11110111000101101111100100001000",
2744 => "00010001000101000000011100010000",
2745 => "00000001000100010000010111111111",
2746 => "00011001111101110000010000000001",
2747 => "00001010000110100000101000001011",
2748 => "00001101000001110000100000000011",
2749 => "00001101000010110000100100000010",
2750 => "00000011000011010000000000000000",
2751 => "11110000000011001111001000001000",
2752 => "00000101000100000000001100000010",
2753 => "00000100111111100000001100000111",
2754 => "00001110000011110000101000000000",
2755 => "00010000000000010001001100010000",
2756 => "00010011000010010000101100000000",
2757 => "00001110000000110000101111111011",
2758 => "11110110111011100001000111111111",
2759 => "00000101111100011111110000000011",
2760 => "11111100000001010000111011110111",
2761 => "11111110111110110000001000010100",
2762 => "11110101111010110000000111111111",
2763 => "00000101111111111110111100011000",
2764 => "11111100000000001111110011111111",
2765 => "00000011111110011111111000001100",
2766 => "00000010111101110000110011111101",
2767 => "00010001000101101111100111111101",
2768 => "00000011000001100001000011111101",
2769 => "11111110000101111111111100010011",
2770 => "00000011111001010000000000000000",
2771 => "00000111111110110000101000101001",
2772 => "00000000111111010000000100000010",
2773 => "11111100111101101111101100011001",
2774 => "11111001000000010000010111111011",
2775 => "11100111000010011111110111111010",
2776 => "11101101111111001110100011110000",
2777 => "00000110000001001111110000000011",
2778 => "11111100111110111111111011110010",
2779 => "00000011111101011111100000001000",
2780 => "00000011111101000000011000000001",
2781 => "00000010111101010000011111100111",
2782 => "11110100111011011111011111110010",
2783 => "11100110111011111111100011110111",
2784 => "11101000111010011110110111101110",
2785 => "11111101111100011111100000000101",
2786 => "11110000111010011111010011110001",
2787 => "11110011111101001110110111111011",
2788 => "11110011111100111111011100000101",
2789 => "11111100111101100000000111110010",
2790 => "11110111111001010000011000000001",
2791 => "11101100111111111111011011110101",
2792 => "00010000111101111111001000010010",
2793 => "11111101111110111111001111111101",
2794 => "00000111111000111111001000001010",
2795 => "11101000111111011111000100000010",
2796 => "11111000000000101110111000000101",
2797 => "11111000111111011111100011110111",
2798 => "11111101000101001111101111111010",
2799 => "11110010000000101111100111111001",
2800 => "00001001000000111111100000001000",
2801 => "00000101111101111111010111111110",
2802 => "00000001000010110000101000000110",
2803 => "00001110111110000000011011111101",
2804 => "00000010111111110000101000000000",
2805 => "11111101111110101111110111111111",
2806 => "11111100000011010000000011111110",
2807 => "11111000111111001111110100000000",
2808 => "00001101000001111111101011111101",
2809 => "00000011000000011111110100000011",
2810 => "11111111000010110000000111111111",
2811 => "00001101111110100000000100000001",
2812 => "00000000000000101111011100000011",
2813 => "11111101000000111111110111111110",
2814 => "11111111000001101111111000000000",
2815 => "11110001111111101111111011111101",
2816 => "00000010111110111111111100000111",
2817 => "00000011111111101111111111111100",
2818 => "11111101111111111111111111111111",
2819 => "00000000111110001111110000000000",
2820 => "11111101111110101110011000000010",
2821 => "11111011111111111111110011110100",
2822 => "11110011000001111111101111111010",
2823 => "11110000111110011111101111111001",
2824 => "11110100111110011111111011111011",
2825 => "00000100111011011111110111111101",
2826 => "00000001000000001111010111111000",
2827 => "11111010111110101111011011110011",
2828 => "11111110111110101111110000000010",
2829 => "11111011111110011111101011110010",
2830 => "00001010111001011111101000000000",
2831 => "00001010000011011111101111111100",
2832 => "00000100111111001111111100000011",
2833 => "11111010000000010000000000001010",
2834 => "11111010111110111111101111111111",
2835 => "11111010000010010000001100000110",
2836 => "11111000000000111111101011111111",
2837 => "00000011000000101111101000011001",
2838 => "11111111111010110000100011111100",
2839 => "00110110111111110000100100000010",
2840 => "00000001000010110010110100000101",
2841 => "00000010000100000000000100010100",
2842 => "11101111111111111111101100000011",
2843 => "11111101000001011111011000010111",
2844 => "11111010111110100000000111111111",
2845 => "00001011111111100000011000100101",
2846 => "00010001111101100000000000001010",
2847 => "11111111000100100000000000000100",
2848 => "00010001000010110001000000001010",
2849 => "11111111000100110000101000001101",
2850 => "00000000111010001111111100001000",
2851 => "00000000000010010001010000010000",
2852 => "11111010000100000000011111111011",
2853 => "00001101000011010000100100001110",
2854 => "00001011111111110000100000000001",
2855 => "00001110000000111111101000000100",
2856 => "11111110000010000001001111111001",
2857 => "00000010000011010000101000001110",
2858 => "00001011111000011111110100000000",
2859 => "11111101000000110000101000001101",
2860 => "00000111000010100000011011110111",
2861 => "00000111000001110000001000001110",
2862 => "00001101111101110000011100000110",
2863 => "00010110111111100000110011111110",
2864 => "11101111000000110010101111101000",
2865 => "00000110000001000000000000001010",
2866 => "00000000111001010000011111110001",
2867 => "00000100111110100000001000010101",
2868 => "11110010000000000000100111111011",
2869 => "00001011111111000000000000010110",
2870 => "00010000111010010000101111111111",
2871 => "00001000000011111111100100000001",
2872 => "11101011000010010001111111101001",
2873 => "00000100000011000000101100011100",
2874 => "00001000110000010000000111101101",
2875 => "00000000000000000000110100011010",
2876 => "00000000000001001111111100000001",
2877 => "00001011000000111111101000010100",
2878 => "00000010111101100000001011111111",
2879 => "00000011000011011111001111111110",
2880 => "11101111000001010000110011101110",
2881 => "11111010000001110000100000000010",
2882 => "00000000111010001111111111110011",
2883 => "00000101111101010000010000000110",
2884 => "11111101000000101111101011111110",
2885 => "00000010111111010000000000000111",
2886 => "00000000111110100000000011111011",
2887 => "11110100000100101110000111111111",
2888 => "11100010111111011110100011011110",
2889 => "00000000000000000000011011111110",
2890 => "11110001111010001111111011111011",
2891 => "00000100111010001111101011101100",
2892 => "11101111000010110000001111111101",
2893 => "00000001111111001111100011110011",
2894 => "11111101111111110000000100000001",
2895 => "11110110111101111111001011111010",
2896 => "11110011111110011111010011110101",
2897 => "00000011111110101111111000001100",
2898 => "00000001111011000000011011111011",
2899 => "00000011111011101111111000000110",
2900 => "11111011111101110000011100000011",
2901 => "11111011000000001111110111111011",
2902 => "11110111111111010000010011111101",
2903 => "11101011111010100000010011110110",
2904 => "11111011111000111111001000000001",
2905 => "11111111111010101111100000000100",
2906 => "00000101111111101111111111111011",
2907 => "11111100111101101111011111110110",
2908 => "11111000111111000000000000000101",
2909 => "11110011111111000000010011101101",
2910 => "11110110111110111111101111111001",
2911 => "11111000111111001111101111110110",
2912 => "00000110111100100000010000000011",
2913 => "00000000111101001111101100000010",
2914 => "11111001111011001111110100000001",
2915 => "11111000111101100000000011111110",
2916 => "00000010111110101111100000000010",
2917 => "11111000111111010000000011111011",
2918 => "11101101000001101111110111111000",
2919 => "11111110111101111111101011111001",
2920 => "00001101111100110000010000001011",
2921 => "11111111111111001111111100000110",
2922 => "11110101000000011111110000000011",
2923 => "11111110000001101111000000001100",
2924 => "00000011111110111110111100000010",
2925 => "11111011000000111111111111111110",
2926 => "00000011111101010000000000000111",
2927 => "11110101111110110000010000000011",
2928 => "11111100000001011111011100000001",
2929 => "11111101000000100000010011101101",
2930 => "00001010000001000000110100000001",
2931 => "00001101111101010000010011101100",
2932 => "11111101000001110001000100000010",
2933 => "00000111000001000000001011111010",
2934 => "11111101111101100000010100000110",
2935 => "00010000111011110000101000000000",
2936 => "11111101111110100001010000000000",
2937 => "00000101111101101111100000000101",
2938 => "11110110000100101111011011111101",
2939 => "11110111111110001111011000000010",
2940 => "00000101111111110000000111111011",
2941 => "11111101111111010000011000010000",
2942 => "00000100110011100000011100001010",
2943 => "00001001111101110001100000000101",
2944 => "11111110000000010000110100000001",
2945 => "11110111000000010000010111111110",
2946 => "00000000111101001111010000000011",
2947 => "11110001000001001111101000000001",
2948 => "11110111000010000000000111111111",
2949 => "00000111000010100000001000001000",
2950 => "00000011111000100000010011111110",
2951 => "00001011000000010000101000000110",
2952 => "00000001000000110001010111111111",
2953 => "00001000000000100000110100010001",
2954 => "11110111111011101111100111111111",
2955 => "11110000000000011111101000001010",
2956 => "00000101000010101111011111110110",
2957 => "00001000000001010000110000010000",
2958 => "00010000111011100000011000000000",
2959 => "00000000000100001111101100000010",
2960 => "11111010111111000001001011110110",
2961 => "00000001000100100000110100001000",
2962 => "00000010111100111111100111111110",
2963 => "11110001111110000000110000001001",
2964 => "00000010000001011111111000000110",
2965 => "00000100000001000000011000001000",
2966 => "00000010111110010000001111111101",
2967 => "11111111000010101111011000000111",
2968 => "00000111111110110000000011111011",
2969 => "00000101000001000000011011111111",
2970 => "00000010111101100000001111110010",
2971 => "00001010000001000000011100000000",
2972 => "00000001000011000000011011111010",
2973 => "00000001000001010000000000000001",
2974 => "00001000111110110000110111111101",
2975 => "00000011000011011110100100000100",
2976 => "11110101111101110000010111101100",
2977 => "00001010000001000000011000010011",
2978 => "00000100111000000000011011100100",
2979 => "00001000111111000000111100001010",
2980 => "11111111000011100000011000000101",
2981 => "00000111000010111111111000000111",
2982 => "00001000000000100000011000000011",
2983 => "00001001000000111111001100001100",
2984 => "11011111111110100001001111100001",
2985 => "11111000000000100000000100001101",
2986 => "11111100111101111111111011011000",
2987 => "00000110000000010000101000010000",
2988 => "11111011000000000000001000000010",
2989 => "11111100000010101111101000010000",
2990 => "00001011111111100000011111111001",
2991 => "11111111000010111101100011111100",
2992 => "11000101111111000000111111010110",
2993 => "11110011000100010000000100000010",
2994 => "11111001111110011111011011001111",
2995 => "11111110111011010000010100010000",
2996 => "11111000111111011111101011111010",
2997 => "00000001111110111111111000010001",
2998 => "00001100111111110000010000000001",
2999 => "11011110000011101100111011110101",
3000 => "11000110000010101110011111011010",
3001 => "11111111000010110000100000001000",
3002 => "00001111000000100000000111001100",
3003 => "00000011111100100000111011111110",
3004 => "00001001111111111111101100000000",
3005 => "00000001111110000000001011101010",
3006 => "11111101000000010000000111101101",
3007 => "11001101000000011101110111110011",
3008 => "00001010111111101100011000001000",
3009 => "11111111111110000000001100001100",
3010 => "11110101000010001111101111010011",
3011 => "11111100111110100000010011101110",
3012 => "11110011000001001111010100000100",
3013 => "00000000111110111111101011011000",
3014 => "11110110111110111111101111111000",
3015 => "11100100111100101111110011110101",
3016 => "11111001111100111111110011111100",
3017 => "11111011111011101111010111111111",
3018 => "11111000111101101111101000001111",
3019 => "11111101111101111111100000000010",
3020 => "00000011111110101110111100000101",
3021 => "11111110111111001111010111110011",
3022 => "11111111111111011111110111110101",
3023 => "11111110111101111111101111111010",
3024 => "00001011111101010000000100010001",
3025 => "00000000111111101111111000000110",
3026 => "11111101111100101111110100000011",
3027 => "11111000000010011111000100000101",
3028 => "00000101111110101110111000000110",
3029 => "11111100111111110000000100000011",
3030 => "00000110000010111111111111110110",
3031 => "11111111000010110000011000000101",
3032 => "11110011000001001111101011110101",
3033 => "00000000000011010000011011111011",
3034 => "00000011111111001110100011110001",
3035 => "11011000000000001111100000000000",
3036 => "00001001111111111111101100000001",
3037 => "00000001111111110001000100000110",
3038 => "11110011111110011111001111110111",
3039 => "00001100111100010010011000000010",
3040 => "11111000111111010000111111110001",
3041 => "00000111111110011111010111111001",
3042 => "11111100000011111111001111111000",
3043 => "11101111111111111110100111111010",
3044 => "11111110111101001111011100000100",
3045 => "11111010111101110000000100000011",
3046 => "11111001110101111111011111111010",
3047 => "00001001111011000001011100000100",
3048 => "11111110000000110000101111111100",
3049 => "11111100111111010000000100001001",
3050 => "11111101000000011111010100000110",
3051 => "11011011111111111110101000000011",
3052 => "00000001111100011111011100001101",
3053 => "11111001111110101111101100001010",
3054 => "11111000111001011111101111111111",
3055 => "00001110000000110000011000000011",
3056 => "11111111000000010000001011111111",
3057 => "00000011111111111111111000000001",
3058 => "00000110111111011111100100001111",
3059 => "11100011000001001111110100000010",
3060 => "00000010000000001111100100001000",
3061 => "11111110000000100000000000010000",
3062 => "00000010111101011111111100000000",
3063 => "00001011000011110000100000000100",
3064 => "00000010111111100000110000000000",
3065 => "00011100000100010000010100001100",
3066 => "11110111111111111111111100001111",
3067 => "11110010000001101111010000001000",
3068 => "11111111000000010000001000001110",
3069 => "00000000000001110000010000001101",
3070 => "00001001000001011111100111111001",
3071 => "00001000000011010000011000000101",
3072 => "00000000111111000001001111111010",
3073 => "00011100000000100000001000010111",
3074 => "00000010000000000000001111101111",
3075 => "11111100000001000001000100001001",
3076 => "11111001000001011111110100000011",
3077 => "00000001000000111111101100001011",
3078 => "00001011000001110000001011101010",
3079 => "00000000111111010000000000000001",
3080 => "11111011111110010000101011110111",
3081 => "00011001000000000000001100001110",
3082 => "00000100000000011111111111000110",
3083 => "00001110000001000000101000001011",
3084 => "11110111000000011111011000001100",
3085 => "00000000000000111111110000000001",
3086 => "00000110000010000000010011101101",
3087 => "11111010111110111110111000000101",
3088 => "00000011111100010000101000001001",
3089 => "00000011111110010000000000000011",
3090 => "11111101111110111110110011001011",
3091 => "00000100111110111111111100001011",
3092 => "11111000000001011110110000010110",
3093 => "11111110000000100000010011111101",
3094 => "00001000000001010000001111101111",
3095 => "11111000000001011101101011111111",
3096 => "00000011111110111111110100000110",
3097 => "11111010111111110000000100000001",
3098 => "00000000111110001110001011100110",
3099 => "00000001111111100000111000001110",
3100 => "00000000000001011110100100000011",
3101 => "11111111000011001111110111111011",
3102 => "00000110000000010000011011111000",
3103 => "11011001000010001101101011111111",
3104 => "11101110111111001100111011110111",
3105 => "11110000111110111111111111100100",
3106 => "00000110111111001110110111011101",
3107 => "11110111111110010000110111101111",
3108 => "00000011000001001110100000000110",
3109 => "11111100000000110000000011011100",
3110 => "11101100000001101111001011110101",
3111 => "11110001110101001110111100000000",
3112 => "00010100111100001100110100011000",
3113 => "00000101111010001111010011110001",
3114 => "11110100000001011111000000000001",
3115 => "11111011111110011110010011010011",
3116 => "11110101111101011111110100000110",
3117 => "11101111111111010000000111010101",
3118 => "11110110111011101110111111101110",
3119 => "11111010111010010000000111111100",
3120 => "00000111111110000000001011111101",
3121 => "00000001111111101111100100000001",
3122 => "11110001111011111111011011111110",
3123 => "11101001111101011110101011110101",
3124 => "11110110111000001110100000000011",
3125 => "11110110111011001111001011111000",
3126 => "11111000111101001111111111111100",
3127 => "00000111111111101110111011111101",
3128 => "00000111111101000000010100001010",
3129 => "00000100111110001111101000000010",
3130 => "11111100111110011110111000000001",
3131 => "11011100000000011111010011111010",
3132 => "00000010111101001110100100000010",
3133 => "11110110000000101111110000000000",
3134 => "11111110000010101111111011110111",
3135 => "00001111111110000000001011111100",
3136 => "11111011111011000000011011111011",
3137 => "00001110111110111111100100000111",
3138 => "11110011000001000000100100000111",
3139 => "00001000000000101111010100000110",
3140 => "11110110111110111111011100000111",
3141 => "11111111111110110000000100010011",
3142 => "11110001110111101111111000000001",
3143 => "00001111111000100001011011111111",
3144 => "11110110111110100000010011110000",
3145 => "00000011111110111111011000000000",
3146 => "11110101000011000000110100011011",
3147 => "11111101111110111110110111111001",
3148 => "11110100111110010000100000010000",
3149 => "11110111111101100000000000000110",
3150 => "11110011110110111110110111111011",
3151 => "00000000111001110000110111110111",
3152 => "11110010111101100000100111110101",
3153 => "00001100111111001111100100000011",
3154 => "11110110111110110001000000000110",
3155 => "11101001111101001110011011111011",
3156 => "11111001111001101111101100010110",
3157 => "11110101111100101111011011111010",
3158 => "11111101110011011111110111110100",
3159 => "11111111111011110000111011111011",
3160 => "11110110111100100000101011110011",
3161 => "00010100111100000000000000010001",
3162 => "11111100111101001110100011101111",
3163 => "11001110111111111111001000000111",
3164 => "00000000111010101110101000010111",
3165 => "11110101111100010000000000000101",
3166 => "11111010111100100000000011110111",
3167 => "00000011000000000000010011111000",
3168 => "11011111111110100000011011011100",
3169 => "00010100111110101111110000001011",
3170 => "11111111000000000000011111110011",
3171 => "11110111111110010000001111111111",
3172 => "11111100111111101110010100010111",
3173 => "11111100111101101111011111111101",
3174 => "11111110111110111111000111110001",
3175 => "00001000111110100000100111110111",
3176 => "11110011111110010000111111110001",
3177 => "00100111000010000000000000010011",
3178 => "11101011111110011111111111110011",
3179 => "11111011111110001111101000001100",
3180 => "11101111111111101110111000010111",
3181 => "11110101111101111111010100001101",
3182 => "11110011000000111111110011110101",
3183 => "11111000111111001111111111111011",
3184 => "00010001111100110000000000000100",
3185 => "00010110111110001111110100000110",
3186 => "11111110000000111111010011100000",
3187 => "11111011000011001111110100000101",
3188 => "11110111111110001110101100010100",
3189 => "00000011111110101111100111111100",
3190 => "11111000000010111111001011110100",
3191 => "11111010111110011111010011111101",
3192 => "00011101111101001111111100001110",
3193 => "11111010000000111111010100000100",
3194 => "11111000000000011111010111101111",
3195 => "11111111000011101111011011111101",
3196 => "11111110111100111110111000000100",
3197 => "11111111111101111111001111111100",
3198 => "00000100000010001111101100001001",
3199 => "11110001111110101110011100000011",
3200 => "00001101111110001111000000011001",
3201 => "11110011111111011111101011111001",
3202 => "00000010000000111110010011110010",
3203 => "11111000000001010000010000000000",
3204 => "00010001000000101111100000000101",
3205 => "11111011000001111111111111110110",
3206 => "00000101000000101111110100000011",
3207 => "11110110000000101110110100001001",
3208 => "00001111111110011110101000011111",
3209 => "00000011111101111111111000000010",
3210 => "00000100000001001110011011110000",
3211 => "11101001000011000000101011111011",
3212 => "00001010000000001110111100000000",
3213 => "11110110000010110000000111100101",
3214 => "11110010111111101111000011110100",
3215 => "11110100111100011111010100000001",
3216 => "00011111111110001110101000011101",
3217 => "11110111111100101111010011110010",
3218 => "00000000000000011110111000010111",
3219 => "11101100000000111110101011100110",
3220 => "00000011111100111110000111111101",
3221 => "11110111111111000000010011101011",
3222 => "11101111111100011111100111110010",
3223 => "11101011111010001111010011101110",
3224 => "00001101111001101110001000000101",
3225 => "00000111110111001111000100000001",
3226 => "11111001111011110000101111110111",
3227 => "11111100000001001110101111101001",
3228 => "11110011111110100000100100000010",
3229 => "11101111000000111111000111101001",
3230 => "11111011111110011111100011111101",
3231 => "00000101111110101111100111111000",
3232 => "11110101111100010000001011111110",
3233 => "00000111111101111111100111111110",
3234 => "11110100111001011111001111110100",
3235 => "11100110111101111110100000000011",
3236 => "11110010111110111111000100000101",
3237 => "11111110111110001111110111111010",
3238 => "11110001110111001111010011110011",
3239 => "00001001111101110000011111110011",
3240 => "11101100111111000000100111101001",
3241 => "00001001111101111111100100000111",
3242 => "11110010111010011111101011111111",
3243 => "11110011111010111110011111111100",
3244 => "11110110111100101111100000000010",
3245 => "11111111111011000000001111111010",
3246 => "11110010110110101110110011101110",
3247 => "00011011110111110010000111101011",
3248 => "11100011111100110001001011100001",
3249 => "00010001111010101111000000001100",
3250 => "11101110000000110010011100010111",
3251 => "11111000111001011110100000000110",
3252 => "11110000111010010000000100001110",
3253 => "11110001111001101111000100010001",
3254 => "11111100110010001110100100000001",
3255 => "00001111111100010001111011110000",
3256 => "11101000111110000001100111100011",
3257 => "00001110111101101110110100000101",
3258 => "11100101111011100010100100100001",
3259 => "00000000111011011110111100001110",
3260 => "11101000111011100000100100010100",
3261 => "11101101111010111111000100010010",
3262 => "11101101101111111110101111111000",
3263 => "00001000111011000001010111101001",
3264 => "11011011111101110000110111011101",
3265 => "00100011111100001110110100000111",
3266 => "11101000111000100010100100010001",
3267 => "00000100111011011110000011111110",
3268 => "11101000111000101111101100010111",
3269 => "11111001111010011110110100001000",
3270 => "11101100110100011111011011111100",
3271 => "00010011111000010001101011101111",
3272 => "11100100111100100001100111100101",
3273 => "00011100111011101110111000000110",
3274 => "11101101111011110010010100011000",
3275 => "00001000111010011110110100000010",
3276 => "11110000111011100000001100010111",
3277 => "11110100111011001110100100001100",
3278 => "11101110111101011110110011111111",
3279 => "00000011111001110000101111101111",
3280 => "11110000111010000000011011110111",
3281 => "00100110111011011110110000000001",
3282 => "11101010111111000001111000010000",
3283 => "00001001111101001110011011111101",
3284 => "11100100111100110001001100010111",
3285 => "11101011111100111111010111111101",
3286 => "11110111111111111111001111110101",
3287 => "00000001111011010000111011110110",
3288 => "00000110111001110000100000001001",
3289 => "00101011111101111111011000000011",
3290 => "11110101000001101111101011111001",
3291 => "11110110000000101111111000000100",
3292 => "11111001111100001111100000011110",
3293 => "11110011111101111111001011110100",
3294 => "11110110000001011111101011111110",
3295 => "11101110111101111111110100000000",
3296 => "00011010111011001110101100010100",
3297 => "00001000111100011111011000000110",
3298 => "11111100000010011110000000000010",
3299 => "11101011000011001111111011111011",
3300 => "11111111111110011111010000000110",
3301 => "11110001000001110000010011101110",
3302 => "00000000000010000000000000000110",
3303 => "11101010000000101110101000001000",
3304 => "00011000111100101110011000100000",
3305 => "11111001111101001111011100000101",
3306 => "00001011000001011101101011110001",
3307 => "11101000000010100000101111111110",
3308 => "00001011000001001111011111111011",
3309 => "11110100000011110000100011101100",
3310 => "11111110000000111111101000001011",
3311 => "11111010111110001111110100000100",
3312 => "00010111111011111111001000100010",
3313 => "00000000111010111111011011101011",
3314 => "00000001000000101111010100001110",
3315 => "11101111000010011111111111101100",
3316 => "00000010111111000000001000001001",
3317 => "11110001000000001111110111110100",
3318 => "11101100111110101111011100001010",
3319 => "00000001111000110000000100000000",
3320 => "00100110110111101111110100101001",
3321 => "11111110111010001111011111111111",
3322 => "00000010111111011111111100100010",
3323 => "11101111000100001110001011111001",
3324 => "11111110111111110000010100001000",
3325 => "11110000111111001111110000000010",
3326 => "11110111111111010000001000001111",
3327 => "11111000111101101111111100000111",
3328 => "00100000000001011111110000011011",
3329 => "00000000111101101111110111111100",
3330 => "00000101000000110000110100001011",
3331 => "00000101000011101111101111111000",
3332 => "00000101000000010000011100000100",
3333 => "11110111000011010000100011110100",
3334 => "11110001111111001111100111111111",
3335 => "11110101111110101111100111111010",
3336 => "11111111111111011110111100000000",
3337 => "11111110111101101111011111110101",
3338 => "11111100111011100000100011111111",
3339 => "00000001111101000000000011111000",
3340 => "11111011111111011110111000000000",
3341 => "11111011000000001111100111110101",
3342 => "11110000111011111111000011111000",
3343 => "11111000111010110000010011101101",
3344 => "11101010111100011111001011101100",
3345 => "00000011111100111111011111110011",
3346 => "11101010111011100001101000001100",
3347 => "00001111111011111111000111100101",
3348 => "11101101111101100001001000000101",
3349 => "11111010111100111110111011110100",
3350 => "11100101110101011111010000001000",
3351 => "00000111111001010001101011110010",
3352 => "11110111111101010000011011110111",
3353 => "11111111111001111111001111111010",
3354 => "11110011111111000010010000101011",
3355 => "11111100111101011110100011110000",
3356 => "11111001111110010001100100010000",
3357 => "11110111111101011110111111111101",
3358 => "11101101101110011110101100001001",
3359 => "00001111110111110001111111110101",
3360 => "11110011111111000000111011110010",
3361 => "00000110111011001110111111111010",
3362 => "11100000111010010010100000100001",
3363 => "00000001111100011101110011111011",
3364 => "11100010111011110001101000001101",
3365 => "11110111111110011110110000000111",
3366 => "11110110101010011111000100001000",
3367 => "00001000111010010001101011111000",
3368 => "11101110000000100000101011101011",
3369 => "11111010111110001110111111011111",
3370 => "11101111110111110001111000100100",
3371 => "11111111111011101110110111110100",
3372 => "11100011111101110001000000010101",
3373 => "11110110111110011110111011111100",
3374 => "11110000110101001111010100000101",
3375 => "00010011111010000001010011110101",
3376 => "11111011111111000000010011110111",
3377 => "11110011111101101111001111001110",
3378 => "11110001111100010001100100011000",
3379 => "00000101111101001110101011110101",
3380 => "11110100111110000001000100001101",
3381 => "11111010111110001111111000001001",
3382 => "11111001111110111111010011111100",
3383 => "00000011000000000000011111111101",
3384 => "11110011111110001111100111110010",
3385 => "00010010111111111111100111100010",
3386 => "11101011111011010001001000000111",
3387 => "00010011111011111110110111101111",
3388 => "11101111111100110000100000010101",
3389 => "11111100111110001111011011111101",
3390 => "11110001000000001111010000000001",
3391 => "11100110111101110000010011110111",
3392 => "00000110111101011110001100000100",
3393 => "00010110111011111111001011100001",
3394 => "11111110000000100001001100000000",
3395 => "11111110000001101111100111100010",
3396 => "00000010111111100000110000011011",
3397 => "11111100111111010000000111011110",
3398 => "11110100111111101111011000001001",
3399 => "11111000111011000000110011111111",
3400 => "00001111111101001110110100010110",
3401 => "11111000111100111111010011010101",
3402 => "11110000000010001111011100001101",
3403 => "11100100000000111111001111101011",
3404 => "11110101111101000000101100011101",
3405 => "11110111111101011111001011110000",
3406 => "11101000000000101110110100001111",
3407 => "11110111111001100000011000000011",
3408 => "00011111111110111110010100011000",
3409 => "11110000111010011111101011010011",
3410 => "00000001000101011110111000010000",
3411 => "11100111000001101111011011100101",
3412 => "00000010111100011111111000001101",
3413 => "11111111111111000000100111110101",
3414 => "11111111111100111110111011111111",
3415 => "00000001111011110000111011111111",
3416 => "00000100111011111111010000000101",
3417 => "11110100111011100000010011010001",
3418 => "11111101000001001111001100001000",
3419 => "11101011111111101111101111110100",
3420 => "11111011111111001111101000001100",
3421 => "00000000111100100000000111111011",
3422 => "11110010111011111110100000001000",
3423 => "00010110111001110010000100000000",
3424 => "00010010000000000000111100001011",
3425 => "11110100111110111111010011101110",
3426 => "11100111000010100000100000100001",
3427 => "11110100111111101101011111111110",
3428 => "11101000111110100000110000000111",
3429 => "11111110111101011110111000001001",
3430 => "00000110111111100000011100010101",
3431 => "00001111000011010000110100010100",
3432 => "00000011000011010000111000000111",
3433 => "00000001000000110000110000000001",
3434 => "00001000000001000000110100011110",
3435 => "00001011000010011111101100001000",
3436 => "00001100000001010001001100000011",
3437 => "00010000000010110000100100001000",
3438 => "00000110111110010000010100001000",
3439 => "11110100000010001111100100000101",
3440 => "00001101000001111111001000001100",
3441 => "11111111000001000000001011111101",
3442 => "00000111111111100000010000001001",
3443 => "11111110000001000000111111111100",
3444 => "11111101000010110000001100000000",
3445 => "00000011000010010000011011110000",
3446 => "11111010000000100000010000000010",
3447 => "11100101111111001111110111111100",
3448 => "11111111000000001101111111111100",
3449 => "11111010111110011111111111101001",
3450 => "00000001000100010000010000010000",
3451 => "00000100111110010000000011110011",
3452 => "00000010000000100000100100000100",
3453 => "11111111111111100000000011101011",
3454 => "00000010111001100000001000001100",
3455 => "11111110111110010000000011111111",
3456 => "00000111000010001111010100001010",
3457 => "11110100111111010000001111101111",
3458 => "00001101111101010000011000010100",
3459 => "11111110000001000000011111110010",
3460 => "00000000000000110001000000000010",
3461 => "11111011000001011111101111110010",
3462 => "11111101110100101111111100001010",
3463 => "00001010111110100001111011110110",
3464 => "11111111000001101111111011111110",
3465 => "11101011000010111111100011000011",
3466 => "11111010111110100000011100101010",
3467 => "11100110111110001111001111101101",
3468 => "11110001111111110001010100000101",
3469 => "00000010111111101111000011111011",
3470 => "00000011110111110000011000001011",
3471 => "11111011000000110000001000000100",
3472 => "00001000000011001110111000001001",
3473 => "11011111000010101111101110110110",
3474 => "00000111111110001111100100100010",
3475 => "11100111111111100000001011101000",
3476 => "00000110000001100001010011111000",
3477 => "00000010000011110000100111110000",
3478 => "11111011111011000000000100001010",
3479 => "11110100000000111111110000001010",
3480 => "00000000000010001110111000000101",
3481 => "11010110000001010000001010110001",
3482 => "00000111111100110000000000011010",
3483 => "11110000000000000000000111100000",
3484 => "00000110000001100000111100000110",
3485 => "00000111000010100000000011110011",
3486 => "11111010000001110000000000001001",
3487 => "00000101000000100000010100000010",
3488 => "00000100000000111111100000000001",
3489 => "00000011111111010000000111010111",
3490 => "11111101111101111111111100010111",
3491 => "00000011111111011111100011111000",
3492 => "00000011000001110000110111111001",
3493 => "00000100000001100000110100000011",
3494 => "11110101000011001111011100000100",
3495 => "11111100111101110001001100000110",
3496 => "00000111000001011110010100000010",
3497 => "11111000111110010000000111000111",
3498 => "00000011000011101110111000001000",
3499 => "11100101111111011110111111100111",
3500 => "00001010111101010001010100010111",
3501 => "00000101111111100000010011110000",
3502 => "11111000111100011111111100001010",
3503 => "11111010111011110000011111111111",
3504 => "00000000111111111110010011111001",
3505 => "11011001111101001111110011001111",
3506 => "11111011000001001111111100011001",
3507 => "11101010111111001110101111101010",
3508 => "11111011111110000000011100001000",
3509 => "00000000111110101111110111110111",
3510 => "11110111111010100000011100000101",
3511 => "00001010111100000001000000000001",
3512 => "00000010000001101111100100000110",
3513 => "11011110111100111111111011101011",
3514 => "11111101111110111111110100011110",
3515 => "11110110000000001111001111111010",
3516 => "11111110111110110000101111111010",
3517 => "00000110111111100000000100000000",
3518 => "11110010111001101111110100000110",
3519 => "00001100111101100001001011111111",
3520 => "11101010000000110000101111011111",
3521 => "00000101111110011111101011110000",
3522 => "11111011111101000001001100010101",
3523 => "00000011111101001110101000000010",
3524 => "11111011111011110001000011111100",
3525 => "00000000111100111111110000010010",
3526 => "11110111111010111111010000001000",
3527 => "00011101111101010010011111111010",
3528 => "00000110000001000010010011101011",
3529 => "00000000000001101111111000000001",
3530 => "11101001111111000001100000010111",
3531 => "11111100000000111110011000010100",
3532 => "11101100111110100001000000001010",
3533 => "11111110111100111111100100011110",
3534 => "00010011111110110001000100011011",
3535 => "00011100000110100001011100001101",
3536 => "00001011001001010010010100001011",
3537 => "00000011000111110001010000000110",
3538 => "00001000000000000001001000100111",
3539 => "00000110000010000000101100100010",
3540 => "00010010000111010000111000000010",
3541 => "00010100000011010000100100100101",
3542 => "00001000000000000000001000001001",
3543 => "00010011000011011111111100001010",
3544 => "00001111000001100000111000010011",
3545 => "00000010000010010000011100010001",
3546 => "00000110111111110000011100010011",
3547 => "00001000000100010000100000010001",
3548 => "00000001000010010000001000000011",
3549 => "00000101000010000000001100011101",
3550 => "00000010111111110000010100001101",
3551 => "00000101000011101111000100000110",
3552 => "00000010000010000000000100001010",
3553 => "11110101000100000000011111111111",
3554 => "11111111000011010000100100001000",
3555 => "00000101000001000000011111111100",
3556 => "00000000000010110001000011111111",
3557 => "00001011000010000000000100000110",
3558 => "00000110000001000000101000001000",
3559 => "11111101000000001110100000001001",
3560 => "00001000000001111110110100000100",
3561 => "11100111000000110000001111110101",
3562 => "00010111000100001111001100000001",
3563 => "11110101000010110000111100000100",
3564 => "00001101000000110000011111111000",
3565 => "00000110000010110000000111101101",
3566 => "00001011000000100000100100000011",
3567 => "11110110000000001111110100000011",
3568 => "00001010000001011110101100001101",
3569 => "11010111000000000000011111010101",
3570 => "00001101000100011110111100011000",
3571 => "11101101000011000000100111101001",
3572 => "00001000000001110000101111101001",
3573 => "00000001000011110000100011101100",
3574 => "00000100000001100001010000000110",
3575 => "00000101000010011111111100001011",
3576 => "00001111000010101111010000010110",
3577 => "11011110000010000000100111010111",
3578 => "00011010000011011110010000000011",
3579 => "11101001000001110001110111110111",
3580 => "00010010000100001111111011110110",
3581 => "00000001000100100000101111111110",
3582 => "00001010000010010000100000000110",
3583 => "00000110000010100000100000000111",
3584 => "00001011000000110000000000001000",
3585 => "11010111000011010000001111010101",
3586 => "00001110000101101110001000010101",
3587 => "11100110000010010000110111111011",
3588 => "00001010000010010000101011100111",
3589 => "00001001000011100001000000000111",
3590 => "11111110111111110000100100010000",
3591 => "00000110111110010001010000000110",
3592 => "00001000000001110000010000000011",
3593 => "11101000000000100000001111010000",
3594 => "00000000000010111111100000011110",
3595 => "11110000000010011111010111110001",
3596 => "00001011000010000000110111111110",
3597 => "00000011000010110001001000000011",
3598 => "00000100111110110000010000001010",
3599 => "00000001111111100000110000000011",
3600 => "00001000000001011111110011111110",
3601 => "11110111111111110000000011011100",
3602 => "11111101000010010000100000100100",
3603 => "11110001000000101111100111110010",
3604 => "00001000111111110000110111111100",
3605 => "00000000000000000000100011111110",
3606 => "00000011111001110000100100000000",
3607 => "00001000111111100000001100000011",
3608 => "11110100000000111111111011111100",
3609 => "11110100111111010000101011101110",
3610 => "00000000111110010000011000001001",
3611 => "11110101111110111111110011111011",
3612 => "00000010111110110001001000001100",
3613 => "11111111000010110000100100000001",
3614 => "11111111111100111111110000000110",
3615 => "00000100111101100000111011110111",
3616 => "11111011000000000000011111101111",
3617 => "00000110111110110000001000000000",
3618 => "00000010111111110000111111111111",
3619 => "00000011000001111111011100000011",
3620 => "00000001111110100000011100000000",
3621 => "00000001111101001111011000000100",
3622 => "11111110111110010000010111111110",
3623 => "00001001000001110000110111111110",
3624 => "11100010000001100001110011010011",
3625 => "00000011000001000000011100001011",
3626 => "11111000111101110001010100011010",
3627 => "00001011111100000000010000010001",
3628 => "11111101000001010000110000001000",
3629 => "00000000111100101111010000001111",
3630 => "11110101111101111111111000001100",
3631 => "00001010111011110000111011111100",
3632 => "11100010000000110001010011011100",
3633 => "00010010111110111111101000001110",
3634 => "11101110111111010001011100110010",
3635 => "00001001111011111110001100001111",
3636 => "11110001111101000001001100000110",
3637 => "11111000111101011111110100010000",
3638 => "00001110111100000001001100010110",
3639 => "00010101000111010001010000010000",
3640 => "00000101000011000001011100000111",
3641 => "11111100000110000000110000010101",
3642 => "00010010111101100000001111111001",
3643 => "11110100000001010001100000010100",
3644 => "00010111000011100000101100000001",
3645 => "00000011000011010001000100010101",
3646 => "00000101111110100000001100010000",
3647 => "11111100000101000000011000000011",
3648 => "00010011000001010000000100010111",
3649 => "00000011000001010000001100001010",
3650 => "00001010111100000000011100010001",
3651 => "11111001000100110000101100000110",
3652 => "00000100000011100000110111111111",
3653 => "00000110000100000000001000000001",
3654 => "00000100000010100000101000001011",
3655 => "11111111000000000000100000001100",
3656 => "00000001000000001111111100000011",
3657 => "11111001111111000000010111111010",
3658 => "00000010000010101111010011111011",
3659 => "11110000000000101111101111111100",
3660 => "00001110000010110000011100000000",
3661 => "00000010000001100000101011111100",
3662 => "00001001000001110000101111111111",
3663 => "11110111000001111111101100000100",
3664 => "00001010111110011111100000001010",
3665 => "11110110000001000000110011110101",
3666 => "00000110000110011101001111111010",
3667 => "11011001000010000000100011111111",
3668 => "00000101000010011111100011110111",
3669 => "00000001000010100000001111110110",
3670 => "00010010000101010000110111111100",
3671 => "11110101000101011111000000001011",
3672 => "00001110000001011111000100010101",
3673 => "11100010000100100000100111101101",
3674 => "00010101000110001101101011110110",
3675 => "11100101000010100010100011111100",
3676 => "00001010000110001110111111110010",
3677 => "00000011000100010000101111110100",
3678 => "00001010000011110000111111111111",
3679 => "11110011000010001111110000001111",
3680 => "00010111000000001111111000010011",
3681 => "11011010000001010000101011101011",
3682 => "00001101000101101101111000000001",
3683 => "11101010000101010001001011110101",
3684 => "00001010000100111111011011110010",
3685 => "00000111000001100000010111110001",
3686 => "00001000000000100000010100000100",
3687 => "00000101000001100001000100001011",
3688 => "00000011000001110000100000000111",
3689 => "11100001111111100000110111100011",
3690 => "11111110000011101110111100001000",
3691 => "11110001000011000000110011110110",
3692 => "00000100000010100000010011110011",
3693 => "00001101111101110000110111111001",
3694 => "00000001111100000000010000000100",
3695 => "00000001000001010000011000001000",
3696 => "11101010111110100000001111111000",
3697 => "11110011000001000000111011101101",
3698 => "11110111000000100000100000001111",
3699 => "11101111111011011111010111111100",
3700 => "11111011000011000000101011111010",
3701 => "00001100111110010000011000000101",
3702 => "11111111111110010000100100001001",
3703 => "00001010000011000000101000000111",
3704 => "11111001000001000001001111111101",
3705 => "11111000000001110000010100000011",
3706 => "00000100000010000001011100001100",
3707 => "00001101000000101111110100001100",
3708 => "00001000000001100001100111101111",
3709 => "00001101000001110000010000001101",
3710 => "00000101111110100000010000000001",
3711 => "00001110000001110000001100000001",
3712 => "11100000000001110001001111011111",
3713 => "00001111000001110000011000011000",
3714 => "11111110111110010010010011110011",
3715 => "00011110000000000000011100010001",
3716 => "11111010000001000001010011111110",
3717 => "00001000000000000000000000010010",
3718 => "11111100111111111111111011110111",
3719 => "00001001000001100000011111111101",
3720 => "11110011000001010001101011011111",
3721 => "00011000000010100000011100100001",
3722 => "11110111111101000010011100001101",
3723 => "00100010000000010000011100010101",
3724 => "00000010000011000001011100000010",
3725 => "00000011111111011111110000010100",
3726 => "11110101000001111111010111111100",
3727 => "00010001000001000000101011110100",
3728 => "11100111000010010001110011011100",
3729 => "00100001000000100000011000110011",
3730 => "11111010111111000010101000010011",
3731 => "00100111111110011111101100010101",
3732 => "00000010111110110001011000000101",
3733 => "11111110111011111111011100011110",
3734 => "11111111111110011111101000001111",
3735 => "00010011000100100001001111111011",
3736 => "11101110000001110001000011100100",
3737 => "00000111000110001111110100000110",
3738 => "11110110111110110001100100001000",
3739 => "00001011111110110000110100001001",
3740 => "11111001111111000001011000000111",
3741 => "00000000111101111111101000010000",
3742 => "00010100111101100001000000000111",
3743 => "00000111000100000000100100000011",
3744 => "11111110000011000001010000000000",
3745 => "00001011000010010000011111111110",
3746 => "00001000000000010001001100001101",
3747 => "11111010000000010001100000010011",
3748 => "00010000000100010010001000000010",
3749 => "00000111000010100000000000010000",
3750 => "00001100111111010000011000001110",
3751 => "00010111000010100001000000010011",
3752 => "00010100000011110001000000011000",
3753 => "00000000000010100000010000010101",
3754 => "00001101111110000000010100000001",
3755 => "00001101000110010001000000011110",
3756 => "00001010000010100001100011111111",
3757 => "00001100000010100000101100011111",
3758 => "00001000000001110000110000000010",
3759 => "00001000000010100000011100000110",
3760 => "00000110000011100000010100000100",
3761 => "11110110000100010000100011111110",
3762 => "00000011001000111110100111110001",
3763 => "11100000000001000000100100000100",
3764 => "00001000000010101111100011111111",
3765 => "00001001000000110000000100001110",
3766 => "00000111000010000000110011111010",
3767 => "11111011000000011111100000000010",
3768 => "00000110000001101111011000001011",
3769 => "11111001000010010000001011111000",
3770 => "00010000001011011101000111101010",
3771 => "11001001000100010000101011111011",
3772 => "00000101111111101110100100000101",
3773 => "00000011000001110000000111111000",
3774 => "00001100000010100000010011111000",
3775 => "11111010000000101111010000001000",
3776 => "00001001111111001111100000001011",
3777 => "11111000000001010000101111111011",
3778 => "00010000000101001100100011011001",
3779 => "11010101000010000000111111111000",
3780 => "00000100000010001101011011111101",
3781 => "00000101000011110000011011111010",
3782 => "00010000000000110001000111110100",
3783 => "11111010111111011111100011111110",
3784 => "00000111111110011111011100000011",
3785 => "00001000000001010000111111111000",
3786 => "00001111000010101110000111101110",
3787 => "11100011000001110001000000000100",
3788 => "00000000000011111110010000001000",
3789 => "00000011000000010000011111111001",
3790 => "00001110111001110000110011111100",
3791 => "00000001111111010000001100000000",
3792 => "11110100111100101111111111111000",
3793 => "11110100111111100000100011111100",
3794 => "00000101000001011110101000000101",
3795 => "11011101000001000000011011111101",
3796 => "11110100000010111110110000000000",
3797 => "00000110000000100000010111111011",
3798 => "00001110111011000000011100000010",
3799 => "11111010000011101111110011111110",
3800 => "11100011111110101111111011101000",
3801 => "11110001000001100000011011110010",
3802 => "00001000111110110001001100000011",
3803 => "11111010111101100000100111111100",
3804 => "11110111000010101111100111111101",
3805 => "00000101000001000000010011111101",
3806 => "00001011111110100000011011111100",
3807 => "00000001000010100000010000000101",
3808 => "11101100111110110000111111101100",
3809 => "00010000000010110000100000001001",
3810 => "00000101000000000000100111101100",
3811 => "00000111111111010000010000001001",
3812 => "11111010000010010000111100000101",
3813 => "11111110111111110000001000000011",
3814 => "00000001000000001111110111110100",
3815 => "00001010000010010000001111111100",
3816 => "11100010000011000001000111011001",
3817 => "00101110000011010000101100100101",
3818 => "00000110111101010001111111110000",
3819 => "00101111111111000000100000010101",
3820 => "11111010000011100000100000000001",
3821 => "00000101111111010000001100001111",
3822 => "00000101000011000000000011100111",
3823 => "00001000000101100000001111110011",
3824 => "11101101000001100001010111011110",
3825 => "00110011000011000000011100100110",
3826 => "11111101111111000010001111111111",
3827 => "00101001111110100000011100011101",
3828 => "11111011000010110000110000000010",
3829 => "00000100111100100000000000010011",
3830 => "11111010000000101111110111111000",
3831 => "00000101000010100000100111110000",
3832 => "11110000000001100000101011101110",
3833 => "00100000000000001111101000100000",
3834 => "00000001111101110010001000001000",
3835 => "00011111111110110000011100001110",
3836 => "11110110111110010000101100001100",
3837 => "11111011111110101111000100001100",
3838 => "00010000111110010000111100000110",
3839 => "00001010000101100000011100000001",
3840 => "11101111001000010001010011110111",
3841 => "00010001000100000000010000010000",
3842 => "11111011111101110010110100001101",
3843 => "00010110111110100001000100011001",
3844 => "11110010000010010010100100000001",
3845 => "00000100000001111111110100010111",
3846 => "00000010000010011111111100000110",
3847 => "00001100000001100000101000000010",
3848 => "00000010000010110000110000000010",
3849 => "00000010000011001111110100000011",
3850 => "11111001000010010000110111111111",
3851 => "00010100000000110000011100001001",
3852 => "11111110000001100000110100000101",
3853 => "00000011000001110000000000000111",
3854 => "00000110000000000000011111101010",
3855 => "00001100111101010001010000000110",
3856 => "11110000111101100000111111111110",
3857 => "00000101000000001111110000001010",
3858 => "00000011000000001111101011110000",
3859 => "11111101111110001111101100001100",
3860 => "00000111111110001110110000000100",
3861 => "11110110111011110000000100001000",
3862 => "00001000000011110000101111101010",
3863 => "11111111111101000000011100000000",
3864 => "11101011111011010000101111110011",
3865 => "00000001000000000000000000000101",
3866 => "00000001000111111111000111100011",
3867 => "11110010111100011111111000000011",
3868 => "00000001111110001110001100000010",
3869 => "11110110111100100000000011111100",
3870 => "00000001000000001111111111110011",
3871 => "00000011000001010000010111111010",
3872 => "11110110111101110000101100000000",
3873 => "00001011111111100000000100001100",
3874 => "00001000000001001111010011101101",
3875 => "11101101111111110001010000000110",
3876 => "11110110111110101101001000000001",
3877 => "00000000111111011111110100000100",
3878 => "00000011111101110000011111110100",
3879 => "00000111111100110000000100000000",
3880 => "11111011111110010001000011111011",
3881 => "00000011000000010000100000001010",
3882 => "00000001000001101110000111101110",
3883 => "11010110000000000001001000001010",
3884 => "11111111000001101101111000000010",
3885 => "00000100111111101111111000001001",
3886 => "00000011110110101111101011101110",
3887 => "00000011000000010000001111110100",
3888 => "11101101111110000000010111101111",
3889 => "00001010000001010000101100000110",
3890 => "00000000111110101111011100011000",
3891 => "11100010111111000000101000000001",
3892 => "11110011000001001101100000000111",
3893 => "00000011111101101111111000000010",
3894 => "00000110110011100000001100000110",
3895 => "00000110111111000000010000000101",
3896 => "11101011000001110000000111110011",
3897 => "11110010000010000000010011111101",
3898 => "11111110111100110000000000000110",
3899 => "11101101111111011111111000000101",
3900 => "11110011000000010000001100000010",
3901 => "00001001111110110000001000000110",
3902 => "00000110110110000000000011111000",
3903 => "00000010000000111111110011111101",
3904 => "11001011111110110000010111010011",
3905 => "00000010000000110000111000000001",
3906 => "11111100111011100000010111111111",
3907 => "11101111111110000000100100000111",
3908 => "11101011000001111111111000000111",
3909 => "00000101111101111111101100001001",
3910 => "00001001111000110000011011101110",
3911 => "00000100000011001111111111110100",
3912 => "11001000111110110000010111001100",
3913 => "00010100000011010000011100000100",
3914 => "00000001111010100010001011110010",
3915 => "00010101111010110000110000001000",
3916 => "11101100000011010000101000001000",
3917 => "00001010111101101111010000000100",
3918 => "00000010000001110000010111111000",
3919 => "00001010000011100000110011101111",
3920 => "11011010000000110001010011011011",
3921 => "00100110000010010000000000010010",
3922 => "00000011111110100011001100000011",
3923 => "00101101111011110000110100001001",
3924 => "11111111000000110001101000000010",
3925 => "00000100111111101111100100001010",
3926 => "00000100000001101111110111110110",
3927 => "00000100000001110000010111110000",
3928 => "11110000000010000000011111110010",
3929 => "00100000000000101111101000001100",
3930 => "11111010111111010011011000010100",
3931 => "00100001111111100000000100001011",
3932 => "11101110000000010001111000000110",
3933 => "11111000111110101111010000001000",
3934 => "11110110111101101111010100000000",
3935 => "11111110000100011111100111111001",
3936 => "11111000000001111111011111110101",
3937 => "00001110000010101111110000000000",
3938 => "00001010111011000001101000001111",
3939 => "00001011111110100000001111110111",
3940 => "00000011111110000001001000000101",
3941 => "11111011111110011111100111111110",
3942 => "11110111111100100000010011111111",
3943 => "11111100000000001111011011111111",
3944 => "11111011000001001111101111111100",
3945 => "00000111000000110000001100001101",
3946 => "11110001111110001111111111111000",
3947 => "00000000111110011111110000000000",
3948 => "11110010000000010000100100000101",
3949 => "11111101000001011111110111111101",
3950 => "11111001000001111111110000000011",
3951 => "00000010111101110000000100000001",
3952 => "00000101111110011111101000000001",
3953 => "00000110111111111111101111111101",
3954 => "00000000000001111111110000001000",
3955 => "00010011000000011111100011111100",
3956 => "11111111111110001111101111111110",
3957 => "11111100111111100000001011111000",
3958 => "11110100000000001111110011111111",
3959 => "11011110000000111111001111110001",
3960 => "11100101111111001110010111101101",
3961 => "11111100111101101111011011110011",
3962 => "11111001111111111111110111111110",
3963 => "00000001111001000000000011101101",
3964 => "00000001111111101110001011111111",
3965 => "00000001111111011111011011100011",
3966 => "11101111111111011110101011101110",
3967 => "11010110111100011110101111101010",
3968 => "11011001111011101101011111100100",
3969 => "11111101111010101111011011100110",
3970 => "11110000111000101111110011111111",
3971 => "00000010110101001110100011011000",
3972 => "11110101111011011101001111111110",
3973 => "11110111111101011111001011001100",
3974 => "11101110110111101110111011101111",
3975 => "11110110111011011111001111111110",
3976 => "11101111111100111111001111110101",
3977 => "00000000111001001111001111111001",
3978 => "11110010110100011111110111100111",
3979 => "11111011111100101101111011111001",
3980 => "11100011110111111110111100000010",
3981 => "11110001111100111111011111110001",
3982 => "11110110110110111111011011101011",
3983 => "11110010111111001111101011110100",
3984 => "11000110111100101111101111100100",
3985 => "00000010111110001111011111111100",
3986 => "11101110111001100000000011100110",
3987 => "11100100110001101110110111110001",
3988 => "11100111111010011100111111111111",
3989 => "11111101111100001111101111110010",
3990 => "00001001110001000000100011100110",
3991 => "11110111111101011111101111101110",
3992 => "11010001111010001111111011100010",
3993 => "00000010111011111111100000000101",
3994 => "11110011111010011111111111100110",
3995 => "11111000110101111111101011111100",
3996 => "11101000111101001101010000000001",
3997 => "11111001111111101111111011111001",
3998 => "00000011110011000000100011101000",
3999 => "11111100111111100000001111111001",
4000 => "10111001111101010000101111010001",
4001 => "11111010000000101111110100000101",
4002 => "11110010111101000000100011100111",
4003 => "11110010110111011111110100001100",
4004 => "11110100000000101101001000000001",
4005 => "00000100111111000000010000000100",
4006 => "11111101101100000000010011101111",
4007 => "00001000000000001111110111111100",
4008 => "11001000111110110000000111011000",
4009 => "11110100000000100000011000001001",
4010 => "11111101110111110000101111011000",
4011 => "11110010111100111111010000001100",
4012 => "11110001111101111101100111111101",
4013 => "11111111000010010000100000000111",
4014 => "00000000110000000000001011101001",
4015 => "00000110000010011111111111110101",
4016 => "10111010111110100000010111000111",
4017 => "11111000000010010000001111111111",
4018 => "11111100111011000000000111010000",
4019 => "11101001110100011111110100001000",
4020 => "11110100111111011100110000000000",
4021 => "00000001111101010000010000000011",
4022 => "11111110111001011111110011101001",
4023 => "11111001000000010000001111101110",
4024 => "11001011111100101111111111011000",
4025 => "11111011000001101111111111111001",
4026 => "11110001111110001111111111110010",
4027 => "11010011110111110000001000000010",
4028 => "11110011111111111100010100000010",
4029 => "00000100111100001111101011111000",
4030 => "11110000111101101110110111101110",
4031 => "11101110111101101111001011110001",
4032 => "11101110111011101111011011110010",
4033 => "11111111111011101111001111110110",
4034 => "11110100111101100000000100000010",
4035 => "11111100111011111111000011111001",
4036 => "11101011111101001110010000000000",
4037 => "11110110111011001111100011110100",
4038 => "00000000111011101111101011111000",
4039 => "11110001111011001111100111111011",
4040 => "11111101000000111111110100000100",
4041 => "00000101111110111111110011111110",
4042 => "11110101111100100000010111111111",
4043 => "00001110111110010000011011111100",
4044 => "11111101111111011110001100000110",
4045 => "11110000111100111111010111111010",
4046 => "11110011111100101111100011111010",
4047 => "11110011111101001111001111111011",
4048 => "00000111111101101111010011111110",
4049 => "11111111111101100000000011110101",
4050 => "11111111111100000000001111110101",
4051 => "11111101111111011111000011111000",
4052 => "11110111111101111110010000000001",
4053 => "11111010111111100000000011110110",
4054 => "00000011000001000000100011111100",
4055 => "00001001000000101111111100000000",
4056 => "00001000111110110000111000000101",
4057 => "00000000111110110000001111111110",
4058 => "00000000000010111111110011111110",
4059 => "11111000111111010000011100001100",
4060 => "00000101000001101110100100000001",
4061 => "00000011000000100000000000001111",
4062 => "00000000000000000000000000000000",
4063 => "00000000000000000000000000000000",
4064 => "00000000000000000000000000000000",
4065 => "11111011000000011111101100000000",
4066 => "11111000000000001111111011111111",
4067 => "00000010111110101111110011111111",
4068 => "11111011111111011111110100000010",
4069 => "11111110000000001111110011111100",
4070 => "11111100111111000000000011111101",
4071 => "11111110000000011110111011111010",
4072 => "00000000111111111111111011111100",
4073 => "00000100000001001111111111111100",
4074 => "11111011000010101111100111111101",
4075 => "11111111000001001111111100000000",
4076 => "11111001000000101111101000000000",
4077 => "11111101111111001111111011111011",
4078 => "00000010111111100000001111111011",
4079 => "00000001111111111110010111111110",
4080 => "11111110111111011111111111111100",
4081 => "00000001000001110000010000000011",
4082 => "11111000000000001111100000000001",
4083 => "00010010000001101111100100001010",
4084 => "11111111000001010000001011111110",
4085 => "00000001111111110000001000000110",
4086 => "00001000111111100000101111111111",
4087 => "11111011000000001111010011111111",
4088 => "00000100000000001111110011111010",
4089 => "11110011000101111111000100000001",
4090 => "11110101111110101111110111111110",
4091 => "00000010111111111111100000000110",
4092 => "11111101111101101111111100000010",
4093 => "00010001111100110000101100001000",
4094 => "00011001111110111111100000000000",
4095 => "00001010111111110001110111111011",
4096 => "11111111111111100000001111110111",
4097 => "00000111111111100000101100000001",
4098 => "11101000000000101111111011111110",
4099 => "00000101000000111111011011111100",
4100 => "11110111000001011111110111111001",
4101 => "11110011000100100000010011111010",
4102 => "00000011111101100000100011101101",
4103 => "11101110000001000000000011111011",
4104 => "00000001000001101110111011100001",
4105 => "11110000111101100000010011111100",
4106 => "11101001111011101111100111111111",
4107 => "11101100111110011111111011110001",
4108 => "11111011111110000000000100000101",
4109 => "00000101111000011111111100000000",
4110 => "00000010111010001111000011110110",
4111 => "11111000111101011111110011111010",
4112 => "11111001111101001111111011110001",
4113 => "00001011111010100000111100000101",
4114 => "11101100111110011111111111111111",
4115 => "00000011111101101110101011111011",
4116 => "11110111000001100000001011111100",
4117 => "11110000110110111111100100000011",
4118 => "11111011111110110000000111101000",
4119 => "11110110000001011111111011111100",
4120 => "00000000000010001111110111101010",
4121 => "11111100111101010000101100000111",
4122 => "11101101111111010000000000000001",
4123 => "00000000111111011110110011111010",
4124 => "11111100111110010000010000000000",
4125 => "00001000111010010000100100000110",
4126 => "00001001111101001111111011101100",
4127 => "00001100000010100000100011111110",
4128 => "00000110000001110001000011100011",
4129 => "00000001111110010000100100001100",
4130 => "11110110111100001111110011111111",
4131 => "11111111111110111111010111110111",
4132 => "11111001111110001111110100000101",
4133 => "11111100111110000000100100000011",
4134 => "00001110111110000000000011111011",
4135 => "00000000000000100000010111111010",
4136 => "11111110000001000000100111110101",
4137 => "11111010000000110000110100010000",
4138 => "11110100111001101111100000000000",
4139 => "11011111111101111111110011101111",
4140 => "11111110111101000000000111111111",
4141 => "00000010111100100000100100001011",
4142 => "00000100111110011110110111111101",
4143 => "00000110000001000000100011111111",
4144 => "11111111000001110001000011111001",
4145 => "11111101000011101111011111110001",
4146 => "11110010111100011111100011111111",
4147 => "11011000111011111111111011100111",
4148 => "11111100111100111111100100000100",
4149 => "11110101000100011111111011101001",
4150 => "00000101111110001110101111111011",
4151 => "11110101111011100000100011111000",
4152 => "11111001111100011111100111111010",
4153 => "11111010110101111111001111100111",
4154 => "11110101111110010000000011111000",
4155 => "11111011111100100000000111111001",
4156 => "11110111111111001111010011111110",
4157 => "11101100110110101110001111110101",
4158 => "11001111111101111110101111111111",
4159 => "11101011111101001100111011111010",
4160 => "11111001111110001111001111111101",
4161 => "11111111111101000000000011111110",
4162 => "11111000000000001111100011111101",
4163 => "00000100111111001111110011111100",
4164 => "11111000111111011111111011111100",
4165 => "11111101111010111111101011111100",
4166 => "11101110111111101111101011111101",
4167 => "11111110111111101101100011111001",
4168 => "11111010111111111111111111111101",
4169 => "00000011000000100000001000000010",
4170 => "00000100000001101111110100000011",
4171 => "00000101000000011111110111111110",
4172 => "11111000000000010000001100000011",
4173 => "11111101000000011111100011110111",
4174 => "00000001000000110000001111111101",
4175 => "11111101000000101110111111111100",
4176 => "00000000111111101111111100001001",
4177 => "00001100111111110000010100001100",
4178 => "00000101000100011111100100000110",
4179 => "11111111000011010000100000000001",
4180 => "11110111000010100000101000001011",
4181 => "00000010111110100000001100000011",
4182 => "00010000000011110000101000010011",
4183 => "00000000000010110000101011111001",
4184 => "00001010000001111111111100010110",
4185 => "00000011000001010000011100000001",
4186 => "00001011000010001111100000001000",
4187 => "00000111000011000000011100000110",
4188 => "11111010000010000000011000000111",
4189 => "00000010000100011111111100000100",
4190 => "00000000000001011111111000010001",
4191 => "00000101111111101111100111111011",
4192 => "00000101000000010000100000000000",
4193 => "00001101000011110000010000000011",
4194 => "00000000000011100000000100000010",
4195 => "11110110000001111111001111110111",
4196 => "11110101000010110000011000000001",
4197 => "00010101000100010000000111110111",
4198 => "00000111111111100000011100000010",
4199 => "00001100000001100000001011111010",
4200 => "11111110000000000000100111111101",
4201 => "00000011111100111111111000000010",
4202 => "00000100000100001110111100000101",
4203 => "00000111000000110000100000000111",
4204 => "11110000111111100000010000001101",
4205 => "11111101111111001111001000000000",
4206 => "11110001000011010000010100010010",
4207 => "11111010000001011111010011110011",
4208 => "00000100000001010000000000001111",
4209 => "00000010000001001111111100000001",
4210 => "00010011000100011110111000000000",
4211 => "11111110000100110001011011111011",
4212 => "11111101000010110000001100011001",
4213 => "00000111111110101111111100000001",
4214 => "00000100000000010000011100010011",
4215 => "00001000111111101111111111110111",
4216 => "00001101111111000000000000011001",
4217 => "00000011000001010000011000001000",
4218 => "00100001000101001111111100000100",
4219 => "11111110000011000010010111111100",
4220 => "11111101000101100000010100101000",
4221 => "11101101111100110000000000000100",
4222 => "00001011000001101111001100100111",
4223 => "00000001000000010000100111110010",
4224 => "00001111000001011111100100100011",
4225 => "00000111111111100000110100000101",
4226 => "00001000000111111111011000001001",
4227 => "11101111000101000001001111110011",
4228 => "11111011000111110000010000010001",
4229 => "00001011111000101111111111111001",
4230 => "00001001000001100000101000011010",
4231 => "00001100000000110000010111111000",
4232 => "00001101000000000000010100010000",
4233 => "00010100000000100000100011111010",
4234 => "11111101000100101101110000000110",
4235 => "11101100000010110000100011100100",
4236 => "00000100000011110000010000001100",
4237 => "00000010111011100000011111100111",
4238 => "00001001000000100000101000010011",
4239 => "11110101111111101111111011111000",
4240 => "00001000111110011111101100001101",
4241 => "00010001000000010000011000000001",
4242 => "11110000000001111101101100000011",
4243 => "11100010000000111110111111010111",
4244 => "11111010000011010000011011111010",
4245 => "00000001111010010000001111101100",
4246 => "00001000111101100000100000001001",
4247 => "00000001000000110000010111111110",
4248 => "00000001111101100000101111110110",
4249 => "11111110111111010000000100000000",
4250 => "11110110111101111111101011111010",
4251 => "11010000111100001110000111100010",
4252 => "11111000111111001111110011111001",
4253 => "11111010111110011111101011101001",
4254 => "11111111111010111111101111101000",
4255 => "11100011111110111111101111111000",
4256 => "00000001111101101110110011110001",
4257 => "11110011000001011111001000001100",
4258 => "11100100111010101111011011110011",
4259 => "11011001110111101110110011100110",
4260 => "11111111111000001111010111111111",
4261 => "11111101111110000000111100000001",
4262 => "00001010111101001110011111110111",
4263 => "00000101111101110001001011111001",
4264 => "11110100111100101111100111101001",
4265 => "11110101111100111111010111100100",
4266 => "11101010111111011111110011110010",
4267 => "11111110110111111111100100000000",
4268 => "11111011111100111111011011111110",
4269 => "11110010110111001111100111111000",
4270 => "11110011111111001111100011111110",
4271 => "11100111111110011111001111111100",
4272 => "11110011111110101110111111110110",
4273 => "00010100000010000000000000000010",
4274 => "11111011000011101111101100000011",
4275 => "11111110000000100000000000000001",
4276 => "11111111000100011111111111111111",
4277 => "11111010000010001111111111111000",
4278 => "11111100000010010000011000000010",
4279 => "11111111111111101111011111111010",
4280 => "00000111000001000000010000000001",
4281 => "11111000111101110000011011111111",
4282 => "00001010000001101111111000000101",
4283 => "00000010000000110000101000000011",
4284 => "11111101000010100000010100000001",
4285 => "11111010111100011111110011111011",
4286 => "11111010111111110000100100001011",
4287 => "00000101000000001111100111111010",
4288 => "00000101111110100000010000000111",
4289 => "11111101111001001111011100000010",
4290 => "00001010000000110000111000000100",
4291 => "00000110000001110000100011111111",
4292 => "11111001000010000000001000001000",
4293 => "00001000000000100000000011111100",
4294 => "11111110000001000000001100001010",
4295 => "11111110000000100000010011111011",
4296 => "00000010000000111111110000001101",
4297 => "00001010111101010000010000000101",
4298 => "00001111000000010000100111111110",
4299 => "00000001000001010001001000000001",
4300 => "11111110000010110000100000001101",
4301 => "00000100000000100000101100000110",
4302 => "00001100000010000001010000001101",
4303 => "11111110000001110000100011111101",
4304 => "00000100000000111111101100010010",
4305 => "11111111110110110000010100000011",
4306 => "00010100111101100000110000000100",
4307 => "00000001000001000001110111111000",
4308 => "00001110000000010000000000100101",
4309 => "00000100111111010000001100001010",
4310 => "00000010111110110000001000001001",
4311 => "11111111000010000000011011111000",
4312 => "00000000000001100000011000010011",
4313 => "00001110111011110000111000000101",
4314 => "00010000000001011111101100000111",
4315 => "11111010000010010010000111110011",
4316 => "00011011000010000000001100101000",
4317 => "00000111111011000000111000001001",
4318 => "00001100000000110000101100011011",
4319 => "11111011000011010000001111101011",
4320 => "00000010000010111111011100010110",
4321 => "00010001111101110000110100000001",
4322 => "00000001000001011110000111111010",
4323 => "11110000000001100000111011111010",
4324 => "00011001000001100000010100101000",
4325 => "00001001110110110000110111111110",
4326 => "00010001111111000000101100010101",
4327 => "11111000000011000000100111100110",
4328 => "00000110000001100000010100001000",
4329 => "00000101000000010000101100000001",
4330 => "11111101000011011110011000000000",
4331 => "11100011000001000000000111101100",
4332 => "00000111000010000000010000011110",
4333 => "00001101111011101111111011100011",
4334 => "00001011000000000001000100001101",
4335 => "00000010000000011111110011111011",
4336 => "00000101000010011111111100000111",
4337 => "00000010000000000000010011110110",
4338 => "11111000000011111101111011111001",
4339 => "11100111111100001111110011010011",
4340 => "11110111000000110000010100000111",
4341 => "11111101111011011111010011010011",
4342 => "00000011111111000000010000000111",
4343 => "11111110000001001111010011111001",
4344 => "00000000111111110000000011111111",
4345 => "00000100111111011111110111111101",
4346 => "11110010000100001101110111111100",
4347 => "11001101111110011110100111011111",
4348 => "11111000000100000000011011111111",
4349 => "00001011111100101111111111010000",
4350 => "00000000111101100000111100000001",
4351 => "00001001000000001111101111110110",
4352 => "00000001000000100000100111111100",
4353 => "00000110000000000000001111110000",
4354 => "11110011000010011101110111111011",
4355 => "10101111111110111110101011000010",
4356 => "11110110000001110000101000001001",
4357 => "00000011111010101111001110111111",
4358 => "11111101111101011111111011111100",
4359 => "11111101111110101111011111111101",
4360 => "00000010000000010000001111111110",
4361 => "00010001000000000000101111110110",
4362 => "11101010000100001111001111111101",
4363 => "11001101000001011101110111011010",
4364 => "11111101000100010000111111111001",
4365 => "00000011111101011111101011001010",
4366 => "00000010111100010000111011101001",
4367 => "00001000000011001111101111110010",
4368 => "00001010000000100000000111101010",
4369 => "11110011000010101111100011101001",
4370 => "11000000111001111110100011111001",
4371 => "11101011110111011101000111110101",
4372 => "11111010110111101111011100000101",
4373 => "11101000000010010000000111101001",
4374 => "00000100111101111110000111101110",
4375 => "11101000111001101111110111111010",
4376 => "11111000111100011111001111010101",
4377 => "11110111000001110000000100000111",
4378 => "00001100111111111111110000000000",
4379 => "00000010000001010000010111111110",
4380 => "11111101111100010000100100000000",
4381 => "00000000000010000000000011111110",
4382 => "00000001000000010000001000000011",
4383 => "11111001000001110000011011111011",
4384 => "00000000000000011111111000001110",
4385 => "00001000111100110000001000000000",
4386 => "00000111000010110000111100000110",
4387 => "00000010111111100000101111111111",
4388 => "00000101000010000000001100000010",
4389 => "00000101000101000000100100000001",
4390 => "00010000000000110000100100000111",
4391 => "11111001111111101111111011111001",
4392 => "00000011111110111111101100000011",
4393 => "00000100110111110000011000001000",
4394 => "00010110000000010001000011111110",
4395 => "11111110111111010001000011111111",
4396 => "00000110000000000000000100000101",
4397 => "00000000000000000000010000001010",
4398 => "11111010000001111111110100001011",
4399 => "00000001000001010000000111111110",
4400 => "11111101000001001111111100010001",
4401 => "00001011110100010000001111111010",
4402 => "00001110111110100001010000000011",
4403 => "11111100111110110001010011111100",
4404 => "11111110111110110000010000001000",
4405 => "11111000111111010000011100001111",
4406 => "11111011111111010000001100000010",
4407 => "11110001000001000000010000000001",
4408 => "11111111111111110000001100001000",
4409 => "00001001110001100000000011111111",
4410 => "00001001111101110001100111111101",
4411 => "11110010111111000001100111110000",
4412 => "11111011111110100000001100010101",
4413 => "00000010111110010000011000010000",
4414 => "11110001000000000000000100000100",
4415 => "00000100111111111111111111111000",
4416 => "11111100111110110000011100000011",
4417 => "00000111101110010000100111111101",
4418 => "00001011111111010000011100000010",
4419 => "11110010111110100001110111110001",
4420 => "11111000000000000000011100010110",
4421 => "11111001110111010001101100010111",
4422 => "00000001111101100000001000001101",
4423 => "11110100000010010000000111110100",
4424 => "11111111000000001111110000001000",
4425 => "00000100110111100000100100001001",
4426 => "00001111000000110000101011111110",
4427 => "11101101000011000000111011110000",
4428 => "11111010000000011111111000000110",
4429 => "11111110111011000001001000000010",
4430 => "00001100000000001111101000001101",
4431 => "00000010111111110000110011010011",
4432 => "00000011111111110000001100010100",
4433 => "00000101111111010000100100000010",
4434 => "00001000000000100000001011111101",
4435 => "11111011000001111111111111110111",
4436 => "11101011000000100000000011111110",
4437 => "00000110111110011111101000001101",
4438 => "11111111111111101111110011111011",
4439 => "00000110111111110000011011011100",
4440 => "11111111000011010000100111111101",
4441 => "00000010000000010000011100000101",
4442 => "11111000000001011111110100000001",
4443 => "11110011000001101111001100000010",
4444 => "11101011111111011111111011101011",
4445 => "11111110000001011111001111111000",
4446 => "11110110111110100000010111111010",
4447 => "00000111000001111111111011100110",
4448 => "00000001000010010000101011110111",
4449 => "00000011000010000000001100000001",
4450 => "11110110000010111111011100000000",
4451 => "11110111000000011110100100000101",
4452 => "11110010000000010000011011011110",
4453 => "00000110111111111110101011011111",
4454 => "11110111000000110000110111101111",
4455 => "00001100000100001110111011110101",
4456 => "00000010000010000000101011110000",
4457 => "00001000000010010000011000000011",
4458 => "11100010000010111101110111111100",
4459 => "00000101111111011101101000010001",
4460 => "11111100111110101111111111101011",
4461 => "00000110111110101110111111100011",
4462 => "00000001000001010000011111100011",
4463 => "11111111000010101110111011111010",
4464 => "00000101000100110000010111011000",
4465 => "00000011000011100000111111101111",
4466 => "11110000111111011111001100000010",
4467 => "11001100111100111110011111110011",
4468 => "00000010111011110000100011101101",
4469 => "00000000000001101111101011100011",
4470 => "00000011111011011111110011101110",
4471 => "00000111000001111111011011111000",
4472 => "11111110111111100000101011101111",
4473 => "11101110111110001110100011011010",
4474 => "11110000111100011111110011101011",
4475 => "11111111110110001110100111111100",
4476 => "11111011111001101110111111111011",
4477 => "11101100111111011101111111111011",
4478 => "11101010111001011101011111101111",
4479 => "11011001110111011011011111111111",
4480 => "11101010111001101110110111100101",
4481 => "00001000111111011111110111111111",
4482 => "11111101000001110000010100000001",
4483 => "00000111000001110000000000000001",
4484 => "00000001000010010000000111111100",
4485 => "11110010111111111111100011111111",
4486 => "11101011000001111111111000000001",
4487 => "11110101000010001111100111111101",
4488 => "00000110000001011111110111111111",
4489 => "11110100000011001111101111111001",
4490 => "00001010111100100000111000000011",
4491 => "11110101000001000000001111110010",
4492 => "11111111111110101111111111111010",
4493 => "11111100000100010000100011110111",
4494 => "00010000111111001111100011111111",
4495 => "00000111111011011111111011111101",
4496 => "11111101111101011111110000000110",
4497 => "11111000110011101111001100000011",
4498 => "00010111111110100001100011111000",
4499 => "11101110000000010000111111110101",
4500 => "00000010111111101111111000001101",
4501 => "11111001111101110000001011111100",
4502 => "11101101111111101111100100000101",
4503 => "11110011111110011111111011111101",
4504 => "00000000111101111111011100010011",
4505 => "11111100110010011111011011111101",
4506 => "00010100111011010001101111111011",
4507 => "11110001111110010000110111110100",
4508 => "00000101111111101111011100001101",
4509 => "11110011000000010000101000100010",
4510 => "11010001111110101110100100000000",
4511 => "11110001111100011111110011111110",
4512 => "11111000111111001111010100001101",
4513 => "11111101110001011111101011111110",
4514 => "00010111111101010001111111111010",
4515 => "11110101111111110001011111111011",
4516 => "11111110000000000000010011111011",
4517 => "11111010111101000000100100111000",
4518 => "11001010111101011111011100000000",
4519 => "11110000111110010000000100001001",
4520 => "00000100111101101111001100001100",
4521 => "11110011101110101111110000000010",
4522 => "00011111111010110010010011110110",
4523 => "00000010111111100001111011111110",
4524 => "11101100111111100000001000000000",
4525 => "11110101111111000000100100101110",
4526 => "11000110111101101110010100000110",
4527 => "11101101111101010000001111111010",
4528 => "00000001111110100000000000010110",
4529 => "11111100110101000000011100001110",
4530 => "00001011111111100001100111111010",
4531 => "11111010000010010000100011111000",
4532 => "11001010000001100000001011100110",
4533 => "00000000000000100000011100101001",
4534 => "11100011111110111111101111111011",
4535 => "00000010000000100001001011101000",
4536 => "00000010000000011111111100000001",
4537 => "11111011111100101111111000001100",
4538 => "00000111111100010001111100000001",
4539 => "11111100000001001111111111111100",
4540 => "11010000111110100000100111101110",
4541 => "11111000000100001111100000100001",
4542 => "11101011111110001111101011111001",
4543 => "11111011111111100001001111011000",
4544 => "00000101000001000000010100000100",
4545 => "11111101111111100000000000010010",
4546 => "00000101111110010000110100000111",
4547 => "11110101000000011111011100000100",
4548 => "11100101111111101111101111010101",
4549 => "00000011000110001111110000100001",
4550 => "11110000111111001111101111110000",
4551 => "00000110111111010001011011010100",
4552 => "00000000000000000000100011111011",
4553 => "00001110000001000000101000000100",
4554 => "11111100000001000000001100001010",
4555 => "00000001000001001110110100001010",
4556 => "11101000000011000000100010111011",
4557 => "00000111000011101110010000000111",
4558 => "11100110000000110000010011101011",
4559 => "00000010000001101111110111111011",
4560 => "11111111000011000000100111101100",
4561 => "00000001000010000000010111110010",
4562 => "11111110111111010000001100000111",
4563 => "00000011111100001110100000000110",
4564 => "11101100000000010000001010111111",
4565 => "00000100000001101100011111110000",
4566 => "11100110000010011111111011100100",
4567 => "00000011000001111101111011110111",
4568 => "00000101000010100000001011101101",
4569 => "11111000000011001111001011100010",
4570 => "11110111111110101111110011110011",
4571 => "11101101110101011110010111110011",
4572 => "11101101111101111111101111011110",
4573 => "00000101000001011101100011011010",
4574 => "11111100111011101110100111101101",
4575 => "00000111111010011100100011110111",
4576 => "11111010111100101111101011110110",
4577 => "11011100110010111110011111101011",
4578 => "10111111110111001110001111101001",
4579 => "00000001110100001011111000000000",
4580 => "11111011101111011101111111111110",
4581 => "11101101110001111101001111111001",
4582 => "10111010111101111101011011001011",
4583 => "11100101110011101011011111111010",
4584 => "11100000111011011110100111000100",
4585 => "11111001000001111111111111110011",
4586 => "00000110111110011111100011111110",
4587 => "11111011111110110000100000000000",
4588 => "11111111111101111111110000000011",
4589 => "11110100000001011111100011110010",
4590 => "11101011111111101111000000000000",
4591 => "11110100111101011110110111111100",
4592 => "11110101111110010000000000001010",
4593 => "11110011000010011111000111110111",
4594 => "00000011111100100001000011110100",
4595 => "11101010111011110000000111101100",
4596 => "11111110111100001110111111111011",
4597 => "11110111000100000001000000001001",
4598 => "00010100111100011111000011110100",
4599 => "00000010111101111111101000000100",
4600 => "11101100111010111111011100000010",
4601 => "11100101110110001110010000000010",
4602 => "00001001110111010001101011101111",
4603 => "11110000000000000000011111110000",
4604 => "11111110111100011110111111111101",
4605 => "11110011000001100001010000100000",
4606 => "11111010111010101110011111110010",
4607 => "11101000111011000001000011111111",
4608 => "11101011111101111111111011111110",
4609 => "11101011110110101110100100000000",
4610 => "00001101110110110010011011110100",
4611 => "00000000111100100000101100000000",
4612 => "00001001111100001111010011111000",
4613 => "11110000000011000000100000100001",
4614 => "11010011111111001101110111110111",
4615 => "11110101111010000000000100001011",
4616 => "11110010111101001110111011111111",
4617 => "11101001101111011111011000000001",
4618 => "00001010111010010010011111110111",
4619 => "00001101111100000000101100001111",
4620 => "11110011111001101110110111110111",
4621 => "11110010000001000000000100110110",
4622 => "11000010000000111110101011110101",
4623 => "11111000111100111111000111111100",
4624 => "11110000111101011111011100000000",
4625 => "11110111101011101111110100010010",
4626 => "00010101111011010010010000000000",
4627 => "00001111000001100001011000010010",
4628 => "11100010111111101111110111111110",
4629 => "11101111111101010000101000111001",
4630 => "11001100000000011111011111111111",
4631 => "11100111000000100000111011110100",
4632 => "11111110111111111111001000001010",
4633 => "11111011101110010000100000010101",
4634 => "00010000111110100001100100001011",
4635 => "00000001000011110000110100000101",
4636 => "11010010000001110000001011101000",
4637 => "00000011111010001111101100110011",
4638 => "11011111000001011111110111111010",
4639 => "11111001000010000001101011100111",
4640 => "00001011000011010000101100001110",
4641 => "00000011111001000000011100001100",
4642 => "00010100000001110010001000010000",
4643 => "11111110000001110000100111110111",
4644 => "11011011000000110000000111101001",
4645 => "11111011111111010000101000101011",
4646 => "11101011111111101111100011111001",
4647 => "11111001111111110001010111100100",
4648 => "00000110111111100000010100010010",
4649 => "00000010111111000000010000010101",
4650 => "00010110000001100010011000000101",
4651 => "11101110000011000001010011110001",
4652 => "11011101000010110000000111011010",
4653 => "11111110000010010001001100101101",
4654 => "00000010111111001111101111111001",
4655 => "00001000000000110001111011100010",
4656 => "00000100000000000000001000001101",
4657 => "00001111111111110000011000001001",
4658 => "00001110000010000001101100001000",
4659 => "11011110000001100000110011101001",
4660 => "11101101000010000000010111001011",
4661 => "11111110000001101111111000001011",
4662 => "11111110111110010000100100000001",
4663 => "11111000000011010001000111110110",
4664 => "00000001000010000000001100000001",
4665 => "00000011111111101111111011101011",
4666 => "00010001111100110001100011111110",
4667 => "10111111111010010000110011000011",
4668 => "00000000111101110000010011011111",
4669 => "11101001000001001110110100000110",
4670 => "11101111111011101110010100000101",
4671 => "11101111111111001111100100000010",
4672 => "11110110111011101111100100001100",
4673 => "00000000111110111111001011110011",
4674 => "00000000111100110000101011110000",
4675 => "11110111111100001111111111111011",
4676 => "11111010111110111111000111101011",
4677 => "11110110000001001101111100010010",
4678 => "11101000111100001111001100000000",
4679 => "11110111111101111101011111111111",
4680 => "11111000111011111111100011111101",
4681 => "11100100110111001110110111110001",
4682 => "10111100111001011110011011111010",
4683 => "11111111111000101100100100000000",
4684 => "11111001111000101111001100000011",
4685 => "11111011110010101111000111101100",
4686 => "11100010111101111111000111010110",
4687 => "11110110110111111110101111111001",
4688 => "11101100111100011111001111010111",
4689 => "11110010000001101111101111111011",
4690 => "11111010000000001111011111111111",
4691 => "11110011000000011111011011101100",
4692 => "11111100111101001111110011111010",
4693 => "00000000111011011111101011111010",
4694 => "00000100111101001111101111110001",
4695 => "11111100111111001111110011111011",
4696 => "11111101111110011111111111111010",
4697 => "11100110111010101110011111111010",
4698 => "11111100111100100001010011110111",
4699 => "11100110000000000000000111101001",
4700 => "00000010111001111110110111110111",
4701 => "11101001111101110001011000000000",
4702 => "00010001111100001110100111110110",
4703 => "11110100111100101111111111111000",
4704 => "11110110111011001111011011111010",
4705 => "11110011111001001110100111110011",
4706 => "00000010111001010000110011101000",
4707 => "11100011111110101111101111100111",
4708 => "00001110111100101110011111111111",
4709 => "11100011000000000001100000000000",
4710 => "00001001111011101110000011110110",
4711 => "11100111111010101111111000001001",
4712 => "11110010111001001110011011111110",
4713 => "11101000000000101110101111110011",
4714 => "00001001111011010000111011101100",
4715 => "11110011000000011111110111110110",
4716 => "00010101111100001111000000000010",
4717 => "11110001000000100000100011111100",
4718 => "11111011111100111110100011111010",
4719 => "11101100111010111111100000000101",
4720 => "11110000111010101111000100001100",
4721 => "11110010111001111111000011111001",
4722 => "00000000111101000000010011111000",
4723 => "00000000111110011111111100000011",
4724 => "00011010111110111111011100000101",
4725 => "11100111000010001111001100001111",
4726 => "11011010000000011110011011111110",
4727 => "11110000111010001111010100001010",
4728 => "11110100111100001111001000000110",
4729 => "11111010101101101111110000001000",
4730 => "00000010111100111111111000000010",
4731 => "00010101000000110000010000011000",
4732 => "00001111111111010000001000001110",
4733 => "11111101111000011111110100011101",
4734 => "11011000000000101111010111111101",
4735 => "11110000111111001111100000000101",
4736 => "11111001111111000000001000000110",
4737 => "00001101110010110000001100001100",
4738 => "00001101000011011111111000000011",
4739 => "00001111000000110001001000000000",
4740 => "11111101000011110000010100010010",
4741 => "00000110111110110000100000011101",
4742 => "11101010000011110001000100001010",
4743 => "00000000000010010000100111100111",
4744 => "00000000000010000000010100001110",
4745 => "00001100111001010000000100000110",
4746 => "00010010000010010001000000001101",
4747 => "11101011000010010001000111100010",
4748 => "11101011000010010000001011110000",
4749 => "11111100111101000001010100011100",
4750 => "11110111111110010000010100001000",
4751 => "11111101000010000001100011011110",
4752 => "00000000000001110000101000001100",
4753 => "00001010000000001111111111111100",
4754 => "00001110000010010001110111111101",
4755 => "11100011111110100001101011011110",
4756 => "11110101000010000000000111111110",
4757 => "00000011000001010001010111110000",
4758 => "00000001111101110000010100001011",
4759 => "00000110111111110000101011101011",
4760 => "00000100111101110000000100010001",
4761 => "00000011111111001111011111101111",
4762 => "00000011000010010000001111111010",
4763 => "11111100111101000001100011101001",
4764 => "00001011111110111111111011111110",
4765 => "00000011111101000000110011111101",
4766 => "11111101111111100000001000010001",
4767 => "00000011000000011111111011110101",
4768 => "11111011000000101111011100000011",
4769 => "11111000111101111111011111110011",
4770 => "11101110111101001111100111101101",
4771 => "11011100111001001111011111010001",
4772 => "00000100111011011111101011100001",
4773 => "11110010111100010000001100000000",
4774 => "11111111111011101110111111110100",
4775 => "11110101111101011111111111111010",
4776 => "11110001111011111111100011110011",
4777 => "11110111111011101111100011111110",
4778 => "11100011111110101110110011111100",
4779 => "11100000111011011110010011100011",
4780 => "11111100111101111111101011110101",
4781 => "11110100111010001111110100000111",
4782 => "11110000111100111111011111100110",
4783 => "11111010000000001111111000000001",
4784 => "11111100111111111111101011101101",
4785 => "11110001111101111111000111110000",
4786 => "11010000111011111110111011110001",
4787 => "00000001110111111101110100000000",
4788 => "11111101111001011111001111111110",
4789 => "11110111111011100000011111101001",
4790 => "11111010111110001111010111101011",
4791 => "11110010111001111111111111111110",
4792 => "11110011111101001111000111100000",
4793 => "00000110000010000000000100000110",
4794 => "00000000000001111111111011111101",
4795 => "00000010000001100000000011111100",
4796 => "11111110000001111111111011110111",
4797 => "00001000111111010000000111111110",
4798 => "00011000000000000000101011110111",
4799 => "00000010000000111111111011111011",
4800 => "00000001111110101111111011111101",
4801 => "11111111111110011111010011111000",
4802 => "11100111111111001111011111111011",
4803 => "11101101000000011110110011110010",
4804 => "11111100111111011111100111101001",
4805 => "11111011111101010000100111110011",
4806 => "00001010111101011111001011110100",
4807 => "11111110111101100000010011111100",
4808 => "00000010111100011111101111101101",
4809 => "11110111111101101111010111101011",
4810 => "11011011111101101101110011100110",
4811 => "11101001111100011110011111100011",
4812 => "00010001111100001111100100000000",
4813 => "11101101111001110000000011101000",
4814 => "00001010111100101110100011111000",
4815 => "11101000111000111110101100000100",
4816 => "11111001111000111110100111101100",
4817 => "11110010111110001111011111101011",
4818 => "11110010111110001110101011101100",
4819 => "11110010111100011111111011101001",
4820 => "00011001111100011111011100011101",
4821 => "11110011110011110000110111100110",
4822 => "00100101111100111110111000000011",
4823 => "11110000111100011111010100001010",
4824 => "11110001111100011111000100000110",
4825 => "11111100110101111111010111101101",
4826 => "11111000000000111111100011101110",
4827 => "11110000111011010000000111110001",
4828 => "00110100111110011111101000100100",
4829 => "11101100110100010001011011101001",
4830 => "00010111111111111111011000000100",
4831 => "11100111111110001111010100010011",
4832 => "11110111111100011111100100000111",
4833 => "11111101110011101111100011110110",
4834 => "11110101111111111110111111110100",
4835 => "00001001111110001111111111111101",
4836 => "00110100000000000000001000011010",
4837 => "11111001111000010000011011110011",
4838 => "11111010000001100000000011111111",
4839 => "11101000000001101111001100010111",
4840 => "11111100000001001111100100000001",
4841 => "00001000110110000000011111111010",
4842 => "00000111000011101111100100000110",
4843 => "11101000111101100001000011100111",
4844 => "00101010000001000000010100100100",
4845 => "00000010111010000000011111111010",
4846 => "11111010000000110000111100001110",
4847 => "11111010000001111111101111110011",
4848 => "00000011111110110000000000001110",
4849 => "00001001111010011111111111110001",
4850 => "00001111000101110001000000000110",
4851 => "11100101000001100001011111011101",
4852 => "11110101000011010000010000001110",
4853 => "11111101111100010000101011110101",
4854 => "11111100111100010000011100010010",
4855 => "11111101111111110000001011101110",
4856 => "00000001000000110000000100001101",
4857 => "00000011111111101111110011111111",
4858 => "00000111000001110000011111111011",
4859 => "11111000000001000001001011110101",
4860 => "00010010000000110000000100001011",
4861 => "11111010111101100001101111110100",
4862 => "00010010111110010000010000010001",
4863 => "11111001000000100000001111110010",
4864 => "00000001000000101111001100001000",
4865 => "11110111000000001111011011111111",
4866 => "11110111111111101111001000000001",
4867 => "11111001111111101111101111111011",
4868 => "00001010111111100000010011110010",
4869 => "00000000111101000000110011001011",
4870 => "00000110000010100000011111111001",
4871 => "00000001111111100000011111111100",
4872 => "00000010111111111111101000000010",
4873 => "00000011111111101111101011111110",
4874 => "11100001000011001110100111111101",
4875 => "11111011000001001110000111110001",
4876 => "11110110111111000000011011100011",
4877 => "00000100111110111111101011011100",
4878 => "00000000000000100000100111100010",
4879 => "00000010000001001111100111110111",
4880 => "00000001111111101111100111100110",
4881 => "00000111000001100000001011110101",
4882 => "11100101000000101110011000000110",
4883 => "11010011000001111100100111111000",
4884 => "00000100000000000000010011101100",
4885 => "00000100111110010000010111011101",
4886 => "00001010111101110000011111011101",
4887 => "11111101000010011111111111111100",
4888 => "00001011000011000000001011011111",
4889 => "11110011000001111111000111100100",
4890 => "11111000111111101111110011110011",
4891 => "00000010111101001110011011111000",
4892 => "00000010000000111111101100000100",
4893 => "11101001000001111111111111100010",
4894 => "00000010111101111101101011100100",
4895 => "11100100111010000000001111111001",
4896 => "11111011111011111111001011101001",
4897 => "00000010111111010000011100001011",
4898 => "11110101000100101111101100000111",
4899 => "00001111000001111111111100001010",
4900 => "11111100000001000000010111111000",
4901 => "00000100000000101110111111110011",
4902 => "11111000000010000000011011111111",
4903 => "00000101000000001111001011111011",
4904 => "00001001000010010000010111110111",
4905 => "00000010000010110000100011111011",
4906 => "11011011000000001110000111111101",
4907 => "11111101111101101110110011110110",
4908 => "00000000111101100000000011110010",
4909 => "11111101111101000000100011111111",
4910 => "00001110111111011111111111110110",
4911 => "00001101000000111110111100000011",
4912 => "11111101111111101111100111100111",
4913 => "11111111111110001111111111111010",
4914 => "11110010000001101101111011101111",
4915 => "11110100111100110000010011110010",
4916 => "00011100111101101111111000011011",
4917 => "11111000111010100001110111110110",
4918 => "00100101000000011111111000000111",
4919 => "11100101111110010000001100000011",
4920 => "00000010111110011110110100001111",
4921 => "11110010111001111111001111111000",
4922 => "11111001111111101110010111110011",
4923 => "11011111000000000000001111100111",
4924 => "00100110111100111111101100011111",
4925 => "11110101110100010001111011101001",
4926 => "00011101111001111111010100000000",
4927 => "11110011111100011111100100010001",
4928 => "11111010111010111111000100000011",
4929 => "11110110110110101111101111110100",
4930 => "11110001111101111111010011110001",
4931 => "11100110111101010000001111011110",
4932 => "00101110111101111111001100100101",
4933 => "11101011110100110010000011100111",
4934 => "00011101111011101111011000000101",
4935 => "11100110111100011111111100010110",
4936 => "11110110111010111111000100000000",
4937 => "11110001110101011111001011110001",
4938 => "00001010111010111111100011110100",
4939 => "00000000111111110001001111111100",
4940 => "00110111111101101111111100111101",
4941 => "11110000110100000010110000000010",
4942 => "00100110000001101111110100010011",
4943 => "11101010111110111111111000000010",
4944 => "11111001111110111111001000010000",
4945 => "00000000110111011111101111110011",
4946 => "00010101000100010000010111111100",
4947 => "11011111111100010010011011011111",
4948 => "00101010000011010000010000011011",
4949 => "11110101110110100010000000000000",
4950 => "00011111111010011111111100010110",
4951 => "11110100111110100000101000001001",
4952 => "00000001111011111111010100010100",
4953 => "11110100111001011111110000000010",
4954 => "00000010000011010000101011111011",
4955 => "00000101111111110001001000000011",
4956 => "00000110000010111111011100010101",
4957 => "11111110111001110001111011111100",
4958 => "00010110000001110000000000001110",
4959 => "11110111111101100000111011110101",
4960 => "11111110111111111111100000001011",
4961 => "00000100111111001111110100000000",
4962 => "11111000000010011111111100001000",
4963 => "00000110111111100000011000001011",
4964 => "00001001000000001111111100001011",
4965 => "00000000111101000000110111111000",
4966 => "00001011000010111111111000001001",
4967 => "11111111000000110000100111101010",
4968 => "00000001000010110000000000000110",
4969 => "00000011000000100000000111111101",
4970 => "11111001000010011110110100000100",
4971 => "11110101111111001111001011111010",
4972 => "00000101000000000000001011101111",
4973 => "00000010111110101110100011100010",
4974 => "11111001000000100000110111111000",
4975 => "00000111000000001111000111110010",
4976 => "00000011000001110000101011111011",
4977 => "00000100000001000000001111111010",
4978 => "11101001000011001110001000000110",
4979 => "00001101111110101101010100001010",
4980 => "00000001000001110000001111110000",
4981 => "00000101111111001110101111011111",
4982 => "11111001000010110000011111100110",
4983 => "00000101000001011111001011110110",
4984 => "00000001000001000000011011011110",
4985 => "00000100000011010000001111100011",
4986 => "11110011000001111111001000000011",
4987 => "11101111111011101110000000000010",
4988 => "11111100000011000000011111101101",
4989 => "00000101000001111111000011011001",
4990 => "11111111111101110000001111100110",
4991 => "00000001000001011111001011111001",
4992 => "11111111111110100000001011101111",
4993 => "11101011111111011111000011101000",
4994 => "11101011111001011111100011110010",
4995 => "11110111110110011110011111111000",
4996 => "11110111110101011111010111111101",
4997 => "11101011000001001110110100000011",
4998 => "11110010111101001110001111110111",
4999 => "11011100111110011101101111111010",
5000 => "11101101111010111111100111100110",
5001 => "00000101000001010000010100000100",
5002 => "00001001111101111111101100001000",
5003 => "00001000111110110000011111111111",
5004 => "00000000000000100000010000001000",
5005 => "11110111000000111111010011110100",
5006 => "00001011000001011111010000001000",
5007 => "11111100111110011111100011111111",
5008 => "11111100111111100000001000000101",
5009 => "11111111111110100000000000000011",
5010 => "00001001000100101111000100001000",
5011 => "00000000000010000000001100000011",
5012 => "11111100000001100000011000000001",
5013 => "11111100111101100000001111111111",
5014 => "00001100000010001111110111111111",
5015 => "11111111000010010000011011111000",
5016 => "00001100000001101111101000000111",
5017 => "11111101111101011111110000000100",
5018 => "00000111111111101111011011111111",
5019 => "00000011000001100000111000000000",
5020 => "00000011000001100000000100001010",
5021 => "00000100111010010001111011111000",
5022 => "00010011000001111111110100001000",
5023 => "11111001111101011111111100000011",
5024 => "00000100111111111111110000001010",
5025 => "11101110111010101111011011111010",
5026 => "11111110111111101110101111110101",
5027 => "11111001111111001111101011110010",
5028 => "00000110111111011111101000001001",
5029 => "00000110110111010000110000000110",
5030 => "00001100111111001111010000000010",
5031 => "00001010111100111111110000001100",
5032 => "11111011111111101111111100000001",
5033 => "11110010111000111111110011111111",
5034 => "00000100111110001111101011110110",
5035 => "11101100111111100000101011101011",
5036 => "00011101111110101111100000011000",
5037 => "11110101110011100001010000000110",
5038 => "00001100111100101111001000000110",
5039 => "00000000111110110000101000001111",
5040 => "11111010111100101111011000001011",
5041 => "11111111110011111111111111110110",
5042 => "00001100111101101111111000000010",
5043 => "11101100111111110001101111101011",
5044 => "00011110111111111111101100011101",
5045 => "11101010110101110001011000010110",
5046 => "00001010111101001111011100010000",
5047 => "11011110000000000000010100000110",
5048 => "11111110111111011111101000010010",
5049 => "11111100110101111111100011111100",
5050 => "00001111000000010000001011111111",
5051 => "11110010111111100001011111111101",
5052 => "00010001000000010000000000000110",
5053 => "11111011110011010000101000001010",
5054 => "11111111111110010000011000000111",
5055 => "11110111000010010001000000001110",
5056 => "11111001000001010000000000010001",
5057 => "11111011111100111111010000000011",
5058 => "00000111000001000001000100000010",
5059 => "00000001000000100001100100000000",
5060 => "00011000000000110000000011111110",
5061 => "11111000111110000000011100000000",
5062 => "11110111000000011111111011111111",
5063 => "11110010111111010000111111110011",
5064 => "00000001111111001111111100010100",
5065 => "00000100000010110000001100000100",
5066 => "11111011000010100000001000001010",
5067 => "00010000111111001111100100001001",
5068 => "11111110000000111111101111101100",
5069 => "00000010000001101111100000010111",
5070 => "11110111000011100000001011110001",
5071 => "00000010000010110000110011101100",
5072 => "00000100000011000000000011110100",
5073 => "00000100000001110000101100000110",
5074 => "11111111111111101111101100000110",
5075 => "00000110111110001110111100001111",
5076 => "11110011111110000000000011100001",
5077 => "00001000000000011111001011111101",
5078 => "11101011000001001111110011101101",
5079 => "00000001000010010000110011110100",
5080 => "00000001000001010000011011110000",
5081 => "00001011000000110001000011111100",
5082 => "11101111000000101111111000010011",
5083 => "00000100000000101110010100001000",
5084 => "11110101000010010000011011011010",
5085 => "00001001000000011110010011110011",
5086 => "11110110000001010000000011101011",
5087 => "00000111000010011110111111110101",
5088 => "00000100000101000000110111101011",
5089 => "11111111000010000000001111110011",
5090 => "11110000111011001110111011111111",
5091 => "11101000111101111110001100000001",
5092 => "00000110111100100000100011101100",
5093 => "00000100000001001111100000001000",
5094 => "11111101111101011111000111101110",
5095 => "00000000111111101111001111111011",
5096 => "11111111000001100000010111101011",
5097 => "11101000111110101110100111101110",
5098 => "11101101111010001111011011110010",
5099 => "11111010110011111101001100000000",
5100 => "11110101111010011111000011111100",
5101 => "11101111111101111111001011101011",
5102 => "11111010111100101101100011011000",
5103 => "11100011111000001101101011111101",
5104 => "11110010111100101111011011100000",
5105 => "00000100000001011111111000000010",
5106 => "11111001000001001111001011111111",
5107 => "00001111111111101111100000000001",
5108 => "11111111000000100000001011111001",
5109 => "11111010111111110000100000000110",
5110 => "00001111000010011111101111111010",
5111 => "11111100000000111111011111111010",
5112 => "00000011111111111111110111111101",
5113 => "00000010000001001111100100000111",
5114 => "11111111000010111111101100000000",
5115 => "11111000000010100000001011111111",
5116 => "00000100000001110000001000000000",
5117 => "11110110111000010001100100000110",
5118 => "00110111111110111111101011111011",
5119 => "11111000000001010000110011110100",
5120 => "00000010000000100000000111111110",
5121 => "00000111111101010000010000001001",
5122 => "00000011000001001111110111111010",
5123 => "00000001000000110000011000000001",
5124 => "00001011000000110000011000001001",
5125 => "00001000110110100010001000000101",
5126 => "00100001000000110000011000001001",
5127 => "00000100000000110000111111111001",
5128 => "00000100000001001111110000001011",
5129 => "00000110111100100000011000000000",
5130 => "00000101000001111111110111111000",
5131 => "11110100000001000000110011110001",
5132 => "11111101000001000000001000001001",
5133 => "00010010110110100010000011110110",
5134 => "00011001111110110000111100001110",
5135 => "00000011000001110000111011111000",
5136 => "00000101111101101111110100001000",
5137 => "00000101110101011111110100001011",
5138 => "00000101000001010000011111111110",
5139 => "11110100000001110000100111101011",
5140 => "11111000111111100000001000000001",
5141 => "11111110110001110001001000011110",
5142 => "00000100111111000000011100000011",
5143 => "11111001000001110000110111101111",
5144 => "00000001000010001111011100001001",
5145 => "11110110110001111111010100001010",
5146 => "00001010111110100000100000001011",
5147 => "11101111000000110000010111110001",
5148 => "11111111111111000000001011101010",
5149 => "11110100110100010000011100011111",
5150 => "11110000111011111111011011110100",
5151 => "11101100000001100001000000000000",
5152 => "00000101000000100000000000001011",
5153 => "11111010110111001111010100001010",
5154 => "00001010111110100000110100001011",
5155 => "00000001000000100000101000000000",
5156 => "00000001111111000000001011100110",
5157 => "11111000111100100000010000100001",
5158 => "11101111000000111111101011111110",
5159 => "11111001111111100001000000001001",
5160 => "11111100000000000000000100000101",
5161 => "00000100111111100000000100001011",
5162 => "00001000111111110001010000000011",
5163 => "00001010111111110000010000000110",
5164 => "11111100111111001111101111011100",
5165 => "11111101000011100000111000101001",
5166 => "11110011000000101111101011111011",
5167 => "00000000000010010000101111110001",
5168 => "11111111000010010000001111111001",
5169 => "00000010111111100000001100001110",
5170 => "11111001111111111111111000000101",
5171 => "00010101000001001111011000010010",
5172 => "11110010111110100000010111001111",
5173 => "00000111000010000000001000100100",
5174 => "11011011000011001111100011101010",
5175 => "00000100000000110000010111110011",
5176 => "00000101000011100001000111110000",
5177 => "00001011111111010000111011111110",
5178 => "00000101111111000000011100001000",
5179 => "11111011000010001111010000000000",
5180 => "11100110000010000000010011000111",
5181 => "00000011000001011110100000001100",
5182 => "11011110000001000000010111101100",
5183 => "00000011000000110000001011111000",
5184 => "00000011000001000000101011110001",
5185 => "00000101111111110000011011110100",
5186 => "11111100111110001111111100000011",
5187 => "11110011111110111111001100000011",
5188 => "11101100111110110000101011010000",
5189 => "11111001000010001100000000000111",
5190 => "11010011111110001111110111101100",
5191 => "11111011000000011110111011111010",
5192 => "00001000000000000000100111101110",
5193 => "11111010000001011111101111111011",
5194 => "11110011111100111110111011111101",
5195 => "00000111110111101110101100000010",
5196 => "11110100111101111111111011110000",
5197 => "00000111000001011110000111110100",
5198 => "11110101111110011110111011110000",
5199 => "00001000111101111101101111111011",
5200 => "11111111111101100000011011101011",
5201 => "11110000000000001111010111110111",
5202 => "11111000111110101111111011110110",
5203 => "00000011111000101111001000000000",
5204 => "11111100111101001111001100000010",
5205 => "11101111111111011111110000000101",
5206 => "11110110111110011110001011111011",
5207 => "11101100111101011111111111111011",
5208 => "11110101111110101111100111101110",
5209 => "00000000000000010000001000010010",
5210 => "00000011000000011111000100000010",
5211 => "00010001000000010000011100000111",
5212 => "11111100000000110000010000000011",
5213 => "00000101000000101111001100000100",
5214 => "11110100000011101111101100001011",
5215 => "11111110000000100000001011111011",
5216 => "00000100000011100000001000000100",
5217 => "11111101111100011111101100001011",
5218 => "00000001111111010000000100000011",
5219 => "00010011000000010000011000001100",
5220 => "11110010000001110000010011111101",
5221 => "00000100111100101111010011111010",
5222 => "11111101000010111111110000000100",
5223 => "00000010000000001111100011111010",
5224 => "00000100000010010000001011111100",
5225 => "00000011111000101111111111111101",
5226 => "00000010000010011111101111111100",
5227 => "00000000111110110000001011111001",
5228 => "11111111111111010000011100000001",
5229 => "00001000111011000001000111111111",
5230 => "00010010111111110000000111111110",
5231 => "11110101111111110000010011111011",
5232 => "00000110111111110000010100000011",
5233 => "00000110110100010000110000001111",
5234 => "00001000000001101111110111111101",
5235 => "11110101000010110000000011111011",
5236 => "00000101000010011111110100000000",
5237 => "00001000111101100010110100100010",
5238 => "00100011111110000000001000000100",
5239 => "11111001000010010010011111110111",
5240 => "00001000000011100000000000001000",
5241 => "00000000110001010000110000010100",
5242 => "00001011000000100000000100001010",
5243 => "00000100000100000000100000000010",
5244 => "00000001000000101111101000000000",
5245 => "11111001111111010010000000101101",
5246 => "00001100000001111111110000001101",
5247 => "11111001111111100010010111101000",
5248 => "00000100000010000000011100001101",
5249 => "00000110110101110000110000001111",
5250 => "00000011000000100000100000001100",
5251 => "00000010000001000000000111111111",
5252 => "11100000000011010000011011100100",
5253 => "11111110000001010001010100111101",
5254 => "11101000111110011111101011111010",
5255 => "11110111000001100010001111111011",
5256 => "00001001000010010000101111111111",
5257 => "00000110111010110000101100010000",
5258 => "00000101111110000000111100000111",
5259 => "00001010000001010000101011111111",
5260 => "11011000000000000000000011100010",
5261 => "11111110000001010000010000111011",
5262 => "11010011111111111111100011111110",
5263 => "11111111000100000001011100000000",
5264 => "00000110000001000001000011111110",
5265 => "00000000111010110000001000010010",
5266 => "00000100111011010000101000000111",
5267 => "00001110000000100000100100001001",
5268 => "11011110111111101111111011100001",
5269 => "11111111000010010000001100101110",
5270 => "11001000000000111111001000000100",
5271 => "11111111111110110001111111111000",
5272 => "00000000000010100000110000001000",
5273 => "00001001111111100000010000000111",
5274 => "11111101111111100000000100001111",
5275 => "00010100000000010000000000001111",
5276 => "11100011000000110000000011100111",
5277 => "00001001000011001110001100011001",
5278 => "11010110000011110000000111111011",
5279 => "00000111000011010000100111110100",
5280 => "00000101000010010000111111111001",
5281 => "11111011000000011111101000010010",
5282 => "00000010111011001111111100000101",
5283 => "00010001111101001111011000000111",
5284 => "11101110000000100000010111100000",
5285 => "00000100000011011110011000011000",
5286 => "11100010000001011111110011111001",
5287 => "00000000000001100000100011111001",
5288 => "00000101000001010000100011111001",
5289 => "11111000111110111111100000000011",
5290 => "00000101111100010000000000000100",
5291 => "11111100111111001111110111111101",
5292 => "11110001111110000000001111110011",
5293 => "11111010000000001111000011110000",
5294 => "11110001111110101111100000001000",
5295 => "11111101111111011111110111111000",
5296 => "11111101111011100000100100000001",
5297 => "00001011000011111111011100000010",
5298 => "00000101000000010000110111111111",
5299 => "00001111111110110000100000000011",
5300 => "11111110111100101111101011111010",
5301 => "00000100000011101111100000000100",
5302 => "00001001000001110000110000000101",
5303 => "00001000111111111110011011111100",
5304 => "00000010111110001111111100001010",
5305 => "11111011111111101111110111111011",
5306 => "11111101111101101111101011111110",
5307 => "00000100000011110000000000000000",
5308 => "11111011000001011111101011111101",
5309 => "11111001111101000000000011111010",
5310 => "00000110111110000000000100000110",
5311 => "11111100000000101110000111111100",
5312 => "11111011111111001111011011111100",
5313 => "00000100000001010000010111111111",
5314 => "00001000000000010000000100000000",
5315 => "00001010000000010000111100001011",
5316 => "00000010000000101111110100001000",
5317 => "11111110000000001111100111111001",
5318 => "00000011111111000000000100000101",
5319 => "11111111111111111110110011111011",
5320 => "11111111111111010000001011110011",
5321 => "00001000111110000000100011111101",
5322 => "00010100111110110000011111111111",
5323 => "00010100111110110001000100010001",
5324 => "00000000111110010000100000001111",
5325 => "00000101000101001111100011111011",
5326 => "11111101000011010000101000001011",
5327 => "00000001000010101111010111110111",
5328 => "00000001000001010000000100010001",
5329 => "11111111111111001111111111111011",
5330 => "00010010000110100000101000000001",
5331 => "00001110000010110000111000001110",
5332 => "11111011000010010000101100000111",
5333 => "00000100000011011111011011111011",
5334 => "00000010000000100000110100010010",
5335 => "00000001000011110000011011111001",
5336 => "00010101111110100000010000001101",
5337 => "00000101110100000000000100000011",
5338 => "00001111000100010000110000001011",
5339 => "00000001000110000000100111111011",
5340 => "11111001000010110000101011111101",
5341 => "00000001111111010000101011011001",
5342 => "00000001000001110000010000001000",
5343 => "00000001111110110001010111110100",
5344 => "00011000111101110000010100001111",
5345 => "00001001111000010000001011111000",
5346 => "00001100000100001111110100001100",
5347 => "11111010001000100000011111110100",
5348 => "11101111000011110001000011111111",
5349 => "00001010111111000000000111100101",
5350 => "00010011000011000001000000001001",
5351 => "11110100000010101110101111101110",
5352 => "00011001000010011111111000001001",
5353 => "11111111111110001111111100010000",
5354 => "00001111000010010000011100001100",
5355 => "11111110001000110000010100000010",
5356 => "11110100000101110000111011110101",
5357 => "00000010111111100000100100000111",
5358 => "11110110000010001111111100000111",
5359 => "11111111000000100000111111101110",
5360 => "00011000111111010000001100001101",
5361 => "00000110000001110000010100000010",
5362 => "00001001111110000000110100000111",
5363 => "11100100001010110000011011101000",
5364 => "11101010000110100000101011101110",
5365 => "11111110000011100000000100001111",
5366 => "11001110111111011111010011111001",
5367 => "00000011111111010001011011110110",
5368 => "00001101111101110000000100000100",
5369 => "00001010111010010000111000001101",
5370 => "00000010111011000000001000000100",
5371 => "11111110000101100000011000000100",
5372 => "11110110000010000000011111111101",
5373 => "11111101111110100001000000000101",
5374 => "11001001000001011111010000000100",
5375 => "11101110000000010001001011111001",
5376 => "00000011000010110000001000001000",
5377 => "00000001000001010000101100000011",
5378 => "00010011000001010001000100001011",
5379 => "00010000000110000000011100010110",
5380 => "11111100000100100000010000000000",
5381 => "00000010000011011111111100001111",
5382 => "11111001000100000000010000001110",
5383 => "11111111000011000010000111110101",
5384 => "00000001000000100000011000010000",
5385 => "00000100111111010000001111111110",
5386 => "00001100000000100000101000000011",
5387 => "11101100000110000000010011111100",
5388 => "11110100000011011111111000000010",
5389 => "11110111000001001110110011111011",
5390 => "11011100111110011111010011111111",
5391 => "11111111111101101111010011111010",
5392 => "00000101111111011111101000000010",
5393 => "00000101000000100000001111111010",
5394 => "00001000000000010000110011110110",
5395 => "11011111111100100000010111101111",
5396 => "11111011111111101111101100001001",
5397 => "11111100000001001111000100000000",
5398 => "11011111111010100000000000000111",
5399 => "11110011000000101110001011110111",
5400 => "11111011111111001111111100000101",
5401 => "11111001000000111111001011111101",
5402 => "00000001111100110000010011110100",
5403 => "00000000111010010000010111111011",
5404 => "11111000111101011111100100000100",
5405 => "11110110000000011111101100000111",
5406 => "11110110111110101111110100000010",
5407 => "11110110111101111110010011111111",
5408 => "11111010111111001111110011111101",
5409 => "11111100111101111111101000000001",
5410 => "11101100111110011111011011111110",
5411 => "00000100000000001110110111111011",
5412 => "11110111111111001111100000000010",
5413 => "11111010111000101111100111110110",
5414 => "11111101000000111111110011111010",
5415 => "11111100111110101110110011111000",
5416 => "11111011000000001111100011110100",
5417 => "00000000000000000000000000000000",
5418 => "00000000000000000000000000000000",
5419 => "00000000000000000000000000000000",
5420 => "11111110000000010000000011111101",
5421 => "00000110000000000000001011111110",
5422 => "11101001111111000000001011110111",
5423 => "11111100000000111111111111111010",
5424 => "00000010111111011111111111110111",
5425 => "11111110111111010000001000000001",
5426 => "00000100111111100000000011111101",
5427 => "11111110111111100000001000000100",
5428 => "00000000111110000000001011111010",
5429 => "00000010111111001111110100000001",
5430 => "11100110111111001111111011111011",
5431 => "11111100111111101111110011111001",
5432 => "00000000111101011111110111111011",
5433 => "11111000111111111111100011111100",
5434 => "11111110000000011111010111111001",
5435 => "00000000000000001111111000000000",
5436 => "11111011111101111111111111110011",
5437 => "00000001111111001111111011111000",
5438 => "11101101111101011111100011110100",
5439 => "11110111111101101111000111111011",
5440 => "11101100111100111111010111110100",
5441 => "11110110111100101110111011110110",
5442 => "11111000111100001110101011110111",
5443 => "11111010111011111111101111110111",
5444 => "11101111111011001111011111101101",
5445 => "00001000111001100000000111110110",
5446 => "11011110111011111111010011101100",
5447 => "11110110111001111111011111111101",
5448 => "11110111111001101110101011101001",
5449 => "11100010111100011110010111110100",
5450 => "11101111111011111110101011111111",
5451 => "11110100111100111111100111111101",
5452 => "11110101111010101110111111100111",
5453 => "00000001111010111111110111100111",
5454 => "11011111111011011111101111100101",
5455 => "11111100111100101110101111111110",
5456 => "11101011111001111110110111101101",
5457 => "11100101111001111110111111110010",
5458 => "11100111111010001110011011111101",
5459 => "11101011111001101110100111111110",
5460 => "11101101111010001110101111110000",
5461 => "11111011111101001111110111100101",
5462 => "11101000111010001111111011110001",
5463 => "11111010111001001110110111110111",
5464 => "11110010111010001111000011101110",
5465 => "11011010111010111111001100000000",
5466 => "11100111111100101110101111111101",
5467 => "11101110111100101110101111110101",
5468 => "11101011111000111110101011101110",
5469 => "11101100110110101111111111101100",
5470 => "11110110111110011111001011110100",
5471 => "11111100111011011111010011110101",
5472 => "11101011111100011111110000000000",
5473 => "11101101111000001110110011101111",
5474 => "11110001111001101111000111111011",
5475 => "11110011111010001110110011101010",
5476 => "11101011111111101110111111110000",
5477 => "11101000110110011111111111101111",
5478 => "11101100111010011110010111110000",
5479 => "00000100111001011110110011110100",
5480 => "11101101111101111111111100000110",
5481 => "00000000111001001111000011100010",
5482 => "11110011111101010000001011111101",
5483 => "11110000111101111111000011100111",
5484 => "11111100111100011110110011110010",
5485 => "11110000111000101111101011101101",
5486 => "11101100111000011111000011101011",
5487 => "11111001111001111111000111110111",
5488 => "11100110110111111111000011111100",
5489 => "11101010111001011110000111101110",
5490 => "11110011111010101111001011111000",
5491 => "11101110111101001111010011110001",
5492 => "11111010111010011111000011111000",
5493 => "11110010111011111111101011110011",
5494 => "11111111111100001111000000000000",
5495 => "11110111111110111111100011111100",
5496 => "00000100110111011111001011111111",
5497 => "11101101111001110000001011110101",
5498 => "11110000000000001111011011111100",
5499 => "11110000111110111110011111111000",
5500 => "11111001111101011111100111111000",
5501 => "11110001111100011111100111111001",
5502 => "11101011111100101111001111101101",
5503 => "11110111111011111111010011111110",
5504 => "11110010111100101111100111110100",
5505 => "11110101111101101111110011111000",
5506 => "11111001000000001111100111111010",
5507 => "11111001111110111111101011110111",
5508 => "11111011111010001111101111110111",
5509 => "11110101111101101111101111111001",
5510 => "11100101111100110000001111111011",
5511 => "11111010111100011111101100000000",
5512 => "11111110111010011110110111110110",
5513 => "11100110111110111111011100000001",
5514 => "11111000111111111110101111111101",
5515 => "11111010111111101111111000000000",
5516 => "11111110111101001111110111111010",
5517 => "00000011000000110000000011111001",
5518 => "11101010111110011111111111111110",
5519 => "11111010111111110000000111111101",
5520 => "11111110111010110000000111111110",
5521 => "11101110111110111111111000000010",
5522 => "11111000000000011111001011111000",
5523 => "11111111111111101111110011111100",
5524 => "00000001111110100000000000000010",
5525 => "11111100000001001111101100000000",
5526 => "11100111111110101111011111111011",
5527 => "11111001000000101111110011111001",
5528 => "00000011111101100000001011111111",
5529 => "00000000111110100000000111111011",
5530 => "11111111000000001111111011111100",
5531 => "00000010111111000000000111110111",
5532 => "11111000111101001111111011110001",
5533 => "11111100111100101111100111111111",
5534 => "11101010111110101111010111110001",
5535 => "11111001111101111111101011111000",
5536 => "00000010111100001111100111101110",
5537 => "11110101111011101111011111110000",
5538 => "00000011111101101111011011111110",
5539 => "00000000111101000000100011110100",
5540 => "00000010111011111111001111111001",
5541 => "11111000111101100000000011110111",
5542 => "11110110111101001110110111111011",
5543 => "11111100111101011111101011101111",
5544 => "11101100111111001111001011111011",
5545 => "11101001111110101111001011101000",
5546 => "11101010111111111110110111111100",
5547 => "11111000111111101111101011110111",
5548 => "11111000111111101111001111110111",
5549 => "11111000111101001111111011111000",
5550 => "11110010111110001110110111110001",
5551 => "00000010111110101111111111101010",
5552 => "11111000111000100000001111110111",
5553 => "11111110111011101111010111011100",
5554 => "11110110111110011111111100000011",
5555 => "11111010111101101111011111110111",
5556 => "11110101000001101110101111101010",
5557 => "11101000111011111111001111101111",
5558 => "11110010111100111111101111101100",
5559 => "00001000111110111110111011110011",
5560 => "11111110111101110000010011110111",
5561 => "00000010111001001111100011101110",
5562 => "11110101111011011111111100000000",
5563 => "11101100111100001111010111101011",
5564 => "11110011111111101110111011101001",
5565 => "11010011111011101110111111110001",
5566 => "11111010111010111101101111110111",
5567 => "00000010111010111111001011111111",
5568 => "00000011111110011110110111110100",
5569 => "11101001111101111111011111111101",
5570 => "11101110111100101110111111111110",
5571 => "11110000111110101111100011011001",
5572 => "11110111000001111110111011111000",
5573 => "11000011000000101111100011111011",
5574 => "00011000111111101100111100010001",
5575 => "00000100111111001111011111110010",
5576 => "00001110000001001111110100001011",
5577 => "11111111000000100000110111101101",
5578 => "00000011111110011111011100000010",
5579 => "11110100111101111111101011010000",
5580 => "11110011000100011111101011111000",
5581 => "11101110111010010000100011111010",
5582 => "00000000111010111101101111111100",
5583 => "11111100111100011111111111101101",
5584 => "00000011000100111111111011111111",
5585 => "00000010111101101111010011100001",
5586 => "00000111111100111111110111111111",
5587 => "11110010111100011111111011010101",
5588 => "11111001000010001110111011110111",
5589 => "11110000000001000000010111110100",
5590 => "00001111111110011111100000010010",
5591 => "00000110111111011111100111101110",
5592 => "11111101000011111111111000001110",
5593 => "11110011000010010000001011110011",
5594 => "11110111000001101111101111111111",
5595 => "11111001111111101111101111110001",
5596 => "00000011111110011111100011111001",
5597 => "11100111111111111111001000000000",
5598 => "00010001111101101111001000010110",
5599 => "11111000111100111111111011110100",
5600 => "00001000000001000000000100000001",
5601 => "11111011000011110000011011101111",
5602 => "00000110000001111111111011111111",
5603 => "11111001000001101111111111101101",
5604 => "11111001111111101111110000000001",
5605 => "11100010111110011110011100000001",
5606 => "00001101000011001110011000000010",
5607 => "11111010000001011111111111110001",
5608 => "11111100000000111111110000000110",
5609 => "11110101000001011111111111101110",
5610 => "11110110000000001111011011111110",
5611 => "00000111000000000000000111101011",
5612 => "00000100111111010000001000000110",
5613 => "11110000000010001111011000000111",
5614 => "00000000000011011110111100000000",
5615 => "00000000000000010000000011111001",
5616 => "00001000111111100000100000000010",
5617 => "00000110000001100000001111110100",
5618 => "00000100000010110000001111111110",
5619 => "00000111000010101111111011110100",
5620 => "11111101000000110000100000001001",
5621 => "00000111111101010000001100000011",
5622 => "11100111000010101111110011101010",
5623 => "11111010000010001111111111111011",
5624 => "11111101000001100000010011110011",
5625 => "00000010111111011111011100000000",
5626 => "00000101000000100000010011110110",
5627 => "00000110111111100000110111111010",
5628 => "11111011111111110000000111110101",
5629 => "00000101111100101111110011111011",
5630 => "11111011111111001111011111110111",
5631 => "11111011111110001111101011111000",
5632 => "00000001111101111111111011111001",
5633 => "11111010111100001111101011110101",
5634 => "00000001111110011111111111111101",
5635 => "11111000111101001111111111111100",
5636 => "00000011111011000000010000000001",
5637 => "11101000111100100000000011111110",
5638 => "11111111111110111111000111111101",
5639 => "11110111111110100000000011110011",
5640 => "11111001111100110000001000000100",
5641 => "11110111111110001111101111110000",
5642 => "11111000000000101111101111111101",
5643 => "11111111111111100000000111101101",
5644 => "11111111000000011111111011111100",
5645 => "11110010111111001111010100000110",
5646 => "11110000000001001111010011110010",
5647 => "11111100111111011111011111110101",
5648 => "11111010111110000000011111110011",
5649 => "00000100111110101111100111111011",
5650 => "11110111111101100000110011110111",
5651 => "11111101111111100000010011110011",
5652 => "00001010000111101111010111110000",
5653 => "11111100000000010000001011111000",
5654 => "11111100000001001111001111111000",
5655 => "00000101111111010000000011111110",
5656 => "11111111000010000000000111110101",
5657 => "00001010111110101111110000000110",
5658 => "00001011111101110000000111111111",
5659 => "11111110111111000000000011111100",
5660 => "11110111001101011110111111101001",
5661 => "11100001111111001110110011110011",
5662 => "00000101111111011110000000000101",
5663 => "00011001000000001111011100001011",
5664 => "00000111001100010000001111111000",
5665 => "00010011111111010000100011111011",
5666 => "00001111111101101111011000000110",
5667 => "11101010111110011111011011101100",
5668 => "11101010001100101111100011101111",
5669 => "11000111111100101101111111101100",
5670 => "00001010111101011101011100001010",
5671 => "00011100111010101111010000100011",
5672 => "00010011001000101111101111101010",
5673 => "00010111000001001111011000000100",
5674 => "00001000111001101110101100001010",
5675 => "11101100111011111111010011101101",
5676 => "11110001001101111111001111101110",
5677 => "11000010111101101101011111110101",
5678 => "00010101111001001011110100010101",
5679 => "00011100111001101111000100011111",
5680 => "00010000001001111110101111101110",
5681 => "00000001000010000000000111101011",
5682 => "00010100111100001110010000001101",
5683 => "11101001111101011111011011010001",
5684 => "11011111000111101110100111101010",
5685 => "11010111111001111111011111110000",
5686 => "00101110111010101100100100101110",
5687 => "00001010110110111110110111110001",
5688 => "00000001001100011110110100000110",
5689 => "11110101000010010000001111001111",
5690 => "00001001111011101110100100010101",
5691 => "11100010111110001111111111011000",
5692 => "11100110000010101110100111110010",
5693 => "11011011111000011110110111110100",
5694 => "00101101111101001100110100101111",
5695 => "00001000110101111111001011110101",
5696 => "00000011000100111111010100001000",
5697 => "11101110000100111111001011100000",
5698 => "00001001111100001111011000000111",
5699 => "11100111111110010000011011011100",
5700 => "11110110000000101110111000000100",
5701 => "11110000111101010000100100000001",
5702 => "00101011111101001101011100110010",
5703 => "11111110111100101111110011100110",
5704 => "00000110000010111111000100011010",
5705 => "11110000000100010000100111011110",
5706 => "00001000000010011111100011111111",
5707 => "11101110000010010000010111100100",
5708 => "11111010000000110000001100000101",
5709 => "00010011111100110001000100000100",
5710 => "00101011000000000000011000101011",
5711 => "11111111000000011111100011111101",
5712 => "11111110000010001111000100010110",
5713 => "11110101000110001111101100000010",
5714 => "00000100000011000000000111111011",
5715 => "11110101000100000000101100001001",
5716 => "00000100000001001111111111111110",
5717 => "00010001111110010001000000000100",
5718 => "00001110000000110001001100001011",
5719 => "11110100000001100000010011111000",
5720 => "00000111000010000000000100001010",
5721 => "00001000111111000000100000001000",
5722 => "00001111000000101111111111111001",
5723 => "11111111000001100000100100001111",
5724 => "00001011000001010000001100000001",
5725 => "00000010000100000000001011111100",
5726 => "00001010111110111111111100000010",
5727 => "00000001000010000000011111111111",
5728 => "11111110000000000000100100001111",
5729 => "00001011111111001111111100001000",
5730 => "11110111000011010000010011110111",
5731 => "00000110000011001111101100000001",
5732 => "00000010111101011111111000000000",
5733 => "11110011000011000000000111111001",
5734 => "11111110111111011111011111111110",
5735 => "11111110111111000000000011111101",
5736 => "00000000111110001111110100000011",
5737 => "11111010111111110000001011111110",
5738 => "11111110000001010000000111111010",
5739 => "00000001000000101111101111110011",
5740 => "11111000111101001111100000000101",
5741 => "00001000111110100000001000001001",
5742 => "00000011000000010000000000000011",
5743 => "11111010000000111111111000001111",
5744 => "11110100111100010000110111111111",
5745 => "11111110000000111111011100001101",
5746 => "11111000111111000000101011111101",
5747 => "00000101111111011111011100001111",
5748 => "00000101000010101111100011111111",
5749 => "00000000000010011110001111110000",
5750 => "11111000000000100000010111110101",
5751 => "11111100000011101111110100000000",
5752 => "11110011111101110000101111111001",
5753 => "00010000111101010000100100001100",
5754 => "00000001000001001111100011111100",
5755 => "11111101000000001110111000000100",
5756 => "00000100001000101111110011110100",
5757 => "11011011000001101110111011111111",
5758 => "00000011000000111110110011111010",
5759 => "00001111000000011111011000001110",
5760 => "00000110000101010000011111110001",
5761 => "00010111000000010000101100000011",
5762 => "00001101111110111111110011111101",
5763 => "11111001111111101111101111101100",
5764 => "11101000001101101111011011111010",
5765 => "11010010111101011101111011110100",
5766 => "00001011111100011101000000001110",
5767 => "00010111111001011111101000010001",
5768 => "00000110001001001111011111110000",
5769 => "00011101000001011111100011111001",
5770 => "00001010111100111110110000000010",
5771 => "11110001000000101110111111011001",
5772 => "11100110001010111111011011110110",
5773 => "11000101110111101100110111110101",
5774 => "00011000000000001011000000010010",
5775 => "00011011111011101111001000001111",
5776 => "00001010000101011110101111110101",
5777 => "00010111111111111111011111011000",
5778 => "00000101111011011110111000000111",
5779 => "11110100111110111110111011001101",
5780 => "11011101001100011111001011111000",
5781 => "11010011110011001101110011110010",
5782 => "00110001111101101001111100101101",
5783 => "11110011110101001110100111101111",
5784 => "00000000000111101101000000000011",
5785 => "00000010000011101110100111000010",
5786 => "00000101111001101101111000000011",
5787 => "11101100111111111111110111000100",
5788 => "11011101001000111110101100000000",
5789 => "11010011110100101110000111111100",
5790 => "00101111111111011010111000110111",
5791 => "11111111111001011111010011010110",
5792 => "11111000000111111101001100000110",
5793 => "11100111000100001110010111001100",
5794 => "11111111111000111110011100000010",
5795 => "11110100111100110000000010111101",
5796 => "11100001000110101110111011111101",
5797 => "11001001111001011110010011111011",
5798 => "00110010000001001001111000110010",
5799 => "11111110111010111111011111001110",
5800 => "11111110000111011110100000010101",
5801 => "11110000000100111111001010100100",
5802 => "00001000111110101111010111111000",
5803 => "11101111111110000000010110111100",
5804 => "11110110000010111111010100000101",
5805 => "11110110111101010000101100000100",
5806 => "00101000000000001100110100101100",
5807 => "11111011111100101111111011100010",
5808 => "11110100000011111111011000010101",
5809 => "11101111000100101111011011001001",
5810 => "11111011111111110000000000000001",
5811 => "11110110111111001111101111011110",
5812 => "11110111000010111111110000000110",
5813 => "00001110111001110001010100001011",
5814 => "00100011111111001111101000100011",
5815 => "00000000111010111111011111101101",
5816 => "11111010000101111111101000100010",
5817 => "11110000000010101111001111110011",
5818 => "00000101111111111111111111111101",
5819 => "11110110111111010000011011111001",
5820 => "00001001111101000000000011111001",
5821 => "00001100000010010000010100000101",
5822 => "00010001111110100000011000011110",
5823 => "11101111000101011111010111110000",
5824 => "00000011111110011111001000010000",
5825 => "11110111000000110000100100001110",
5826 => "11111001000001001111101011111101",
5827 => "11111001000001001111111000001101",
5828 => "00001001111101101111101100001010",
5829 => "00001010000101000000011000000100",
5830 => "11101000000010111111111100000110",
5831 => "11110100000011111111111011111001",
5832 => "11111101111111100000010011101001",
5833 => "11111000000001000000010100000100",
5834 => "00000100000001001111110011110100",
5835 => "00000110000000000000100000000110",
5836 => "11111110111110001111101011111111",
5837 => "11110011000001000000000011111001",
5838 => "00000111000000001111011000000111",
5839 => "11110111111111101111111100000001",
5840 => "00000000111011100000010100000000",
5841 => "11111010000010011111111100001011",
5842 => "11111100111101101111011111111110",
5843 => "11111101000000001111100111110111",
5844 => "11110110000001011111100011110001",
5845 => "00000000111111101111010011111101",
5846 => "11111011111110100000110111111101",
5847 => "11111010111110111111100100000010",
5848 => "11101100000001011111101011110011",
5849 => "00001000000000001111000011111111",
5850 => "11111101111011011110001111111001",
5851 => "11111000111101111111010000000101",
5852 => "00000010000011101111111100000000",
5853 => "11101101000001101101100000000010",
5854 => "11111110000001000000000000000101",
5855 => "11111111111110111111110100000110",
5856 => "11110100111110100001000111111111",
5857 => "00001111000000010000011100001101",
5858 => "11110011000001101111011100000000",
5859 => "11111101000001001111100011111110",
5860 => "11111110001000100000000000000011",
5861 => "11100101000001011101011111111101",
5862 => "00001010000000001110000100001110",
5863 => "00000010111110101111110000000000",
5864 => "11111011000010000000110011111111",
5865 => "00011110111111100000110111110100",
5866 => "00000110000001010000011111111110",
5867 => "11111110000001011111111111101111",
5868 => "11101100001011001111100100000011",
5869 => "11010111111010001110001011111100",
5870 => "00011010000000001100010100010110",
5871 => "00000100111011111111110111111010",
5872 => "00000110000111110000000000000011",
5873 => "00011011000010101111111111011100",
5874 => "00000010111110000000010011110110",
5875 => "11110111000010101111100111011100",
5876 => "11101110001000011111011100000010",
5877 => "11101110111001011110111100000011",
5878 => "00011100111111001100111100011110",
5879 => "11110100111100001111101011101010",
5880 => "00000111000100001110010100010111",
5881 => "00000100000011000000000011011101",
5882 => "00001000000000000000010011110101",
5883 => "11110011000001110000000011110000",
5884 => "11100101000110111110110111111111",
5885 => "11101101110101100000010011111110",
5886 => "00100010111100001101010000100011",
5887 => "11100001111010011110111111101010",
5888 => "11110111000101001101110000000101",
5889 => "11110111000011001110010111100000",
5890 => "11111001111000111111000100000010",
5891 => "11110110111101101111011011100001",
5892 => "11111000000111011111011100000101",
5893 => "11100110111101011111010111111111",
5894 => "00100011111111001101110100100010",
5895 => "11100011111100111111010111101111",
5896 => "11111100000110011101010011111111",
5897 => "11101101000010101111101011101001",
5898 => "00000011111110011110110011111001",
5899 => "11111001111110001111110111100101",
5900 => "11111011000110001111110000000101",
5901 => "11011101111101111110011111111100",
5902 => "00100001111111111100011100011110",
5903 => "11010111111101110000001111010110",
5904 => "00010001000101001101011000001000",
5905 => "11110011000010000000000111011100",
5906 => "00001110000001001111010011110010",
5907 => "00000001000010000000001111011010",
5908 => "11101110000001111111001000001010",
5909 => "11101111111010101111111011111111",
5910 => "00100100111111111101111000100001",
5911 => "00001001111100011111110011101101",
5912 => "11111100000010101110111000010000",
5913 => "11101011000011001110111111101010",
5914 => "11111110111100100000000111111011",
5915 => "11111101111111001111111011101001",
5916 => "11110111000000001111100000000001",
5917 => "00000100111000110000110000000000",
5918 => "00001000000000001111110000001110",
5919 => "11110111111100011111001111101001",
5920 => "11111001000010111111011100011100",
5921 => "11110111111111101111001111111000",
5922 => "00001011111101110000010011110111",
5923 => "11111101111110001111101100000011",
5924 => "00000100111100000000000100001011",
5925 => "00001000111101000000010100000000",
5926 => "11110111111111110000100000001111",
5927 => "11111011000000101111010000010101",
5928 => "11110101111110101111100100001001",
5929 => "11110011111110010000001000001000",
5930 => "11110000111111001111110000000010",
5931 => "11110100111111011111010100001010",
5932 => "00001011111100100000000011110011",
5933 => "00000001000001111111111111110100",
5934 => "11100001111110000000011011111101",
5935 => "11111010000000010000010111111010",
5936 => "11110101111110101111101111111011",
5937 => "11100010111101100000010000010010",
5938 => "11110100000010011111001011111100",
5939 => "11111100111110101111100100001010",
5940 => "11101101000000011111001011110011",
5941 => "00001011111010000000101111110110",
5942 => "11111111111110000000000011111101",
5943 => "11110111111100011111100000001001",
5944 => "11111110000001001111101111110011",
5945 => "11111000000000101111010100001010",
5946 => "00000000111100011111111011111010",
5947 => "11110001111111001111111000000110",
5948 => "11111001000010001111000000001000",
5949 => "11111011000001000000001100000000",
5950 => "00001011111111111111110100001100",
5951 => "11111001000000011111100100000100",
5952 => "11110000000011011111101100010110",
5953 => "11111001000011011111110100000001",
5954 => "11101011000001000000010011111010",
5955 => "00000000000010101111011011111111",
5956 => "11111101111011011111111000000010",
5957 => "11100000111111111101100000000111",
5958 => "00001000111111001110011000001111",
5959 => "11111000000000010000011011110101",
5960 => "11111101110111110000100100000100",
5961 => "11110000111111100000000111111000",
5962 => "11110011000000110000011111111010",
5963 => "00001011000001110000001111100110",
5964 => "00001010000100100000101000000000",
5965 => "11110111000001101101111100000110",
5966 => "00001001000001001111010100001110",
5967 => "11111111000001000000100111110111",
5968 => "00000010000001011111001111111011",
5969 => "11101111000000100000110011110000",
5970 => "11111100000101000000001111101100",
5971 => "00001010000010000000101011110010",
5972 => "00010001000110100000111100000111",
5973 => "11111000000001111111100000001000",
5974 => "00000100000001011111011100001000",
5975 => "11101011000010000000011111100010",
5976 => "00000100000011011111000000000001",
5977 => "00000001000001010001001011110001",
5978 => "00000001000100100001010011110010",
5979 => "00000100000001110000010111111011",
5980 => "11111110000111100000001100001001",
5981 => "00000100111110110000011000000100",
5982 => "00010110111111011110011100011000",
5983 => "11101110000000010000011011011001",
5984 => "00000001000100011111001100000100",
5985 => "00000110000101101111111011100000",
5986 => "00001111000000110001000011101001",
5987 => "00000100000000100000011111110011",
5988 => "11110010000011111111110111111101",
5989 => "11101010111101011111001111111000",
5990 => "11111001111111111110000011111100",
5991 => "11101101111100101111011011100100",
5992 => "11110100000011100000110000000000",
5993 => "00001110111110111110111011101101",
5994 => "11111010111110000000010011111111",
5995 => "00000011111101101111011111100000",
5996 => "11110110000010000000011011111100",
5997 => "11010010000001001101101000000011",
5998 => "00001110000010011100101100001110",
5999 => "11101010111111100000001011111001",
6000 => "00000110000000101110010011100000",
6001 => "00000001000001110000011011110001",
6002 => "11111101111110111110111011111010",
6003 => "00000011111110101111101011011110",
6004 => "11111010000101110000011100000011",
6005 => "11100000111101111101010000000101",
6006 => "00100110000000111101000000011111",
6007 => "11011111111100110000001100001100",
6008 => "00001101000011011110000111111001",
6009 => "00000001000010010000100111101110",
6010 => "00001000000001011111100011101101",
6011 => "00000000000001011111110011101110",
6012 => "11111000000010011111111011111110",
6013 => "11110001111100101111001111111111",
6014 => "00011110000010011110100100100000",
6015 => "11100100111101111111111011110111",
6016 => "00000100000011001111101100011011",
6017 => "11110101000001110000000111101110",
6018 => "11111110000001011111110011111011",
6019 => "11111111000001101111111111111000",
6020 => "11110011111111101111110100000101",
6021 => "11110111111011101111110011111101",
6022 => "11111011000000111110110100001011",
6023 => "11111100111110001111010111100011",
6024 => "11111001000000010000111100011001",
6025 => "11111111111110001110101011101001",
6026 => "00000101111101000000101011111011",
6027 => "11111010111100001111011011110011",
6028 => "11110000111100101111010011111101",
6029 => "11110100111100111111001011110100",
6030 => "11110111000000001111001111101011",
6031 => "00000111111101111111001111110001",
6032 => "11101110111100110000101111111000",
6033 => "11111101111110101110010011111101",
6034 => "11110101111100100000100011111110",
6035 => "11111000111100001111000011111010",
6036 => "11101011111011111111000011110110",
6037 => "11110001111111111111011011110111",
6038 => "11101011000000001110111111110111",
6039 => "11111101111111101111001011111011",
6040 => "11110010111001101111100111111111",
6041 => "11101100111110101110101011110101",
6042 => "11101101111011111111001011111001",
6043 => "11110110111101101111010111110100",
6044 => "11111000000000101111100111111001",
6045 => "11110011111111000000011111111001",
6046 => "00000001111111101111100000000001",
6047 => "11111110111110011111011011111011",
6048 => "11110111000010110000011100001011",
6049 => "00000010111100111111100011110111",
6050 => "11111110111110011111110111111000",
6051 => "11111000111110011111101011110110",
6052 => "00000111111011000000100000001110",
6053 => "11101001000100101101011100000110",
6054 => "00001011000010001110111000010000",
6055 => "11111011000010010000101000000000",
6056 => "00000010111001101111100100000011",
6057 => "11110000000011000000101111111111",
6058 => "11110010000011000001101011111011",
6059 => "00001010000011100000001011110010",
6060 => "00001111111010110000110100000001",
6061 => "00000001000110101101011100000110",
6062 => "00000001000011100000000100000011",
6063 => "11111011000010100001011011111101",
6064 => "00001010111000101110011111111001",
6065 => "11100000111111100000011100000001",
6066 => "11110110000100011111100111110010",
6067 => "00001110000000110000001100001110",
6068 => "00010000000010010000100100001100",
6069 => "00000100000101011110111100001001",
6070 => "00001000000000111111011000000100",
6071 => "11100011000011010000110011111001",
6072 => "00001011111111011110000000001101",
6073 => "11100110000010010000110011111011",
6074 => "00001111000011110000100011101000",
6075 => "00001000000001110000100100000111",
6076 => "00000111000011000000010100001000",
6077 => "00001010000001000000001000001111",
6078 => "11110011000001001111101011110110",
6079 => "11111011000011110000101011101110",
6080 => "00000000000000101101011100000000",
6081 => "11101110111110101111110111110111",
6082 => "00000001000010010000010011011001",
6083 => "00001101000001100000111000000101",
6084 => "00000101000010000000100100001000",
6085 => "00010001000010110000111000001001",
6086 => "11011110000001100000001111011110",
6087 => "11111000000000100000110000000111",
6088 => "11111111111110011111110000000111",
6089 => "00000110111111101111110000000111",
6090 => "00000110000011100000101011110111",
6091 => "00001101111101100000010000001100",
6092 => "00001010111111100000101000000000",
6093 => "00000001000011111111101011111001",
6094 => "11011011000010000000001011100000",
6095 => "00010011000011010000001100000111",
6096 => "11111010111011110000010011100110",
6097 => "00001111111001110000001000001101",
6098 => "11101100000000111111111000000101",
6099 => "00000110000000111111101000000100",
6100 => "11111111111101110000111011111011",
6101 => "11100000000000101100011111111010",
6102 => "11111111000011001101100100000010",
6103 => "11110011000001110000110011101101",
6104 => "00001001111001111110101111011101",
6105 => "11111101000001000000101111110001",
6106 => "11111101000010111111010011101111",
6107 => "00001000000010000000001111010101",
6108 => "11111001000010100000110100000011",
6109 => "11111100111100011111100100000110",
6110 => "00010101000100111111011000010110",
6111 => "11100001111110100000010011111110",
6112 => "00010100000010101111100111110001",
6113 => "00001011000011000000011011110010",
6114 => "00001101111111110000000011011111",
6115 => "00001001000001110000010111110111",
6116 => "11111000000000110000011000000111",
6117 => "00010010111111000000110100000110",
6118 => "00011000000010010000111100001111",
6119 => "11110101000001101111110100000111",
6120 => "11111110000001100000001100001101",
6121 => "00001001000001101111110000001111",
6122 => "00000111111111000000001111101011",
6123 => "00000010111110011111111100011001",
6124 => "11111110111111000000010100001000",
6125 => "00010100000000100001010011111101",
6126 => "11110110000011110001010111110111",
6127 => "11111011000001001111111100000111",
6128 => "11110100000000100000010000010001",
6129 => "00001100111110001111011000010000",
6130 => "11110100111111000000001000000100",
6131 => "11111111111110101111110100011001",
6132 => "11111001000000101111010100000001",
6133 => "00010010111110000000111011111001",
6134 => "11101001000000000001000111101001",
6135 => "00000011111111011110101100010001",
6136 => "11101010111111110001000000000000",
6137 => "00001011111101101111010000010010",
6138 => "11110001111010100000010011111100",
6139 => "11111010111101111111011100010110",
6140 => "11110100111010001111100111111010",
6141 => "11111111000010000000000111111000",
6142 => "00001101000001011111100100000111",
6143 => "11111101000000101111100000000001",
6144 => "00000000111000011111101111110101",
6145 => "11110010111111110000001011111100",
6146 => "11111010000000001111011111111111",
6147 => "11110101111111111111110111111010",
6148 => "11110111111111011111110000000010",
6149 => "00001110111110001111101111111100",
6150 => "00010010111111010000010100010000",
6151 => "11111110111110001111110100001001",
6152 => "11111000111111000000000000000111",
6153 => "00000000000011001111001100001100",
6154 => "00000101111111010000101111111100",
6155 => "00000000000000100000001000010100",
6156 => "00010010111000110000111000000001",
6157 => "00010100000100011111101000001101",
6158 => "11111100000010100001011000000010",
6159 => "11111010000110010000111000001110",
6160 => "00010011110110100000000011110011",
6161 => "11111000111111010001110000001100",
6162 => "11111110000001100000000011110010",
6163 => "00001010000001000000010100010010",
6164 => "00010000111000110000111100000000",
6165 => "00001011000100110000010011111111",
6166 => "11110110000001000000111111111000",
6167 => "11111011000101000000101100001000",
6168 => "00001000111001101110100011110111",
6169 => "11101010111111000000011100001101",
6170 => "11111110000011111111011111110010",
6171 => "00000111000001100001000000001010",
6172 => "00001101111100100000111100000100",
6173 => "00001000000010010000011000001101",
6174 => "11111000111111110000101011111001",
6175 => "11101010000001110000110100000000",
6176 => "00010001111111001110011111111010",
6177 => "11110100000000010000101100000001",
6178 => "00010000000010100000011111100101",
6179 => "00001000111111110001010100010010",
6180 => "00001011111111001111111000000011",
6181 => "00001110000001100000100000000100",
6182 => "11011000111111000000010011011101",
6183 => "11101111000010100000101011110011",
6184 => "11110111111110011111101111101011",
6185 => "11111100111011001111010000000101",
6186 => "11111001000001000000000011011110",
6187 => "00001001111110010000100100000111",
6188 => "00000110111011010000100100000011",
6189 => "00010100000010100000010011111010",
6190 => "11011111000000000000110011011111",
6191 => "11100000111111110000100000010110",
6192 => "11111101111011110000011011110010",
6193 => "00001001111100111111011000001101",
6194 => "00001000111111011111110111111110",
6195 => "00000111111111100000010100010000",
6196 => "00000101111100001111111000000101",
6197 => "00010001000001110001000111111100",
6198 => "11111011000000110001011011111000",
6199 => "11101100000010010000000000001101",
6200 => "11111101111110100001000011110000",
6201 => "00010110000001011111111000011000",
6202 => "00000000000001110000100011101110",
6203 => "00001001000000111111111100011101",
6204 => "00001011111001110000010100001000",
6205 => "00010000000000010000000000001001",
6206 => "00010001000000110000100000000001",
6207 => "10111111000011010000000111110100",
6208 => "00000111111100001111010011110000",
6209 => "11101000000001110000001100001010",
6210 => "00000000000000100000001011110100",
6211 => "00000101000001110000001100001001",
6212 => "00000100111111100000110100000011",
6213 => "00001000111111000000100000000010",
6214 => "00000100000000100000100011111100",
6215 => "11001111000001010000110011101010",
6216 => "00000110000000011111000100010110",
6217 => "11111000000001000000001000001000",
6218 => "00001010000001101111001111011010",
6219 => "00000111111111110000011100000101",
6220 => "11111011111110110000000000001101",
6221 => "00001000111101100000100000000001",
6222 => "00000000000010110000011111110110",
6223 => "11101001000010010000001011110001",
6224 => "11111101000001000000110100011001",
6225 => "00001001000000001111000000000000",
6226 => "00001000111110100000010111101110",
6227 => "00000111111111011111011100000011",
6228 => "11111100000000001111111100000101",
6229 => "11111011111011100000000111111101",
6230 => "11111000000010010000000111111111",
6231 => "00000100111110101111110111111100",
6232 => "11110111000010010000000100010101",
6233 => "00001100111110011111000111111011",
6234 => "11111011111101010000011100000111",
6235 => "11111010000000101111100011111010",
6236 => "11111001111111001111000011111010",
6237 => "11111111111111001111101111101100",
6238 => "11100101111101111111100111100101",
6239 => "00001011111110001111100000000111",
6240 => "11110111111101100000111011111111",
6241 => "00001011111101001111110100000011",
6242 => "11101110111101110000011011111111",
6243 => "11111111111101111111000111111010",
6244 => "11111110111011101111101011111011",
6245 => "11110101111111111111111111111101",
6246 => "00000011111101100000001000001010",
6247 => "11111011111101011111010011111110",
6248 => "11111100111011001111100111110101",
6249 => "11101111000000100000110000000001",
6250 => "11111000111101010000010011111001",
6251 => "11101111111110111111100111111001",
6252 => "00000011111101111111110011111011",
6253 => "00001111111111010000011111111100",
6254 => "00001101111110110001010100010011",
6255 => "11111110111111111111101100001010",
6256 => "00000001111011100000001100000101",
6257 => "11110011000000110000001000000000",
6258 => "11111101111111110000000111111110",
6259 => "11111001111101111111111000000001",
6260 => "00001100111001010000001111111001",
6261 => "00001111111110100001100011111111",
6262 => "11111110111110000001010011111000",
6263 => "11111111000000000000000000000011",
6264 => "11111010000000010001000100001100",
6265 => "00000100111111110000001100000111",
6266 => "11111111000001010000010011110111",
6267 => "11111000000001000000100100001001",
6268 => "00001001111001100000100000000010",
6269 => "00001000000001010000111000000101",
6270 => "11111011000000100000101111111001",
6271 => "11111001000011010000001100000110",
6272 => "00000000111111101111101100000101",
6273 => "11101110111101110000001000000110",
6274 => "11111000000000110001011111110101",
6275 => "00000110000001110000101000000100",
6276 => "00000000111001110000010011111010",
6277 => "00000011000000010000100000000000",
6278 => "11101001111111000000101111110011",
6279 => "11111000111111010000011000000011",
6280 => "00000100111101011110001011011111",
6281 => "11100101111111111111010100000000",
6282 => "00000010111111111111011011111010",
6283 => "00000101111101110000101000000100",
6284 => "11111100111010001111110100000011",
6285 => "11111110111111000000010111111011",
6286 => "11110001111110101111100011101110",
6287 => "11110001000000110000000011101111",
6288 => "11101110111001101111011111110101",
6289 => "11101111111100101110101011111000",
6290 => "11101110111100101111100011111101",
6291 => "00000010111110111111111011111001",
6292 => "00000101111100000000100100000001",
6293 => "00000100000001010000010111111110",
6294 => "11110000000000000000100111110001",
6295 => "11111001000010000000011111111111",
6296 => "11111001111001110000010011101010",
6297 => "00010010111101101111010000000011",
6298 => "00001000111101100000001100000100",
6299 => "00000111111110100000011000000101",
6300 => "00001001111010010000011100001001",
6301 => "00000101000000100000100100000100",
6302 => "11110110000000000001001011111111",
6303 => "11110010111111010000010100000101",
6304 => "00000010000000110000111111101111",
6305 => "00001110111110000000000000001101",
6306 => "00000000000001010000110100000100",
6307 => "00000100000000110000000100000110",
6308 => "00000100111110110000100100000000",
6309 => "00001000000000110000110000001100",
6310 => "00000010000010000000110111111101",
6311 => "11101000000000100000010011110111",
6312 => "00000010000000011111011011101110",
6313 => "11111111000000100000011100001110",
6314 => "00000100000001100000010100000111",
6315 => "00000001000010100000011000001000",
6316 => "00001001111111010000100000000101",
6317 => "00001011000000010000011011111110",
6318 => "11111100000001011111110111111000",
6319 => "11010011111111110000011111110110",
6320 => "00000110111110000000000011111101",
6321 => "11111100111111100000000100000111",
6322 => "11110111111111001111011111110110",
6323 => "00001010111110011111110100000011",
6324 => "00000011111110100000001100001101",
6325 => "00010110111111100000100000000010",
6326 => "11110010000010100000111111110101",
6327 => "11101011000010110000000000000001",
6328 => "11111010111111000000001100001011",
6329 => "00000101111110001110110100001100",
6330 => "11110110111110011111110111110110",
6331 => "11111111111101111111110000011001",
6332 => "11110100000000111111100100001100",
6333 => "00000101111101110000001111111011",
6334 => "11111000111111110000100000000100",
6335 => "11101110000000101111011100000010",
6336 => "00001000000000111111110100000111",
6337 => "00000011111101111111000100001001",
6338 => "00001110111011101111111111111000",
6339 => "11111000111111010000100100001010",
6340 => "11111101111101001111100000001000",
6341 => "00001001000000000000010111110111",
6342 => "11101110111111110000000000000001",
6343 => "11111110111110111111001011111110",
6344 => "11110001111111110000001000000001",
6345 => "00000011111110001111010011111110",
6346 => "11111101111010011111111011111101",
6347 => "11111010111101011111100100000111",
6348 => "11111000111100101111011111110011",
6349 => "11111100111100010000010111101101",
6350 => "11110101000000111111010111111111",
6351 => "11111110111110011111011111111000",
6352 => "11101100111110010000000000001000",
6353 => "11110011111101001111110011111011",
6354 => "11100001000000100000000111111110",
6355 => "11110101111101101111001111111010",
6356 => "11111011111101011111101100000001",
6357 => "00001101111111000000000111111010",
6358 => "11111101111111110000100100000000",
6359 => "11111001000000011111111100000010",
6360 => "11111110111001111111110011111010",
6361 => "11110100000000101111110100000101",
6362 => "11111110111111010000100111111011",
6363 => "11111101111111101111110000001001",
6364 => "11111101000000011111101111110110",
6365 => "11111110111110110000001111110110",
6366 => "11111111111111000000000011111100",
6367 => "11111100111111001111111100000100",
6368 => "11110010000011000000110000000010",
6369 => "11100000111110001111010111111111",
6370 => "11110100111110111111100011111010",
6371 => "11111110111101011111010011111011",
6372 => "11111011111010111111011111110110",
6373 => "00000101111111000000101000000100",
6374 => "00000011111110000000010000000011",
6375 => "00000001111111101111100100000111",
6376 => "11111001111111110000100000000100",
6377 => "11100010000000011111001000000001",
6378 => "11101110111111101111110111111010",
6379 => "11111110111110110000000100000001",
6380 => "11111101110111101111100100000010",
6381 => "00000111111110100000111011111011",
6382 => "11111001111110101111111011111011",
6383 => "11111000111110001111110011101110",
6384 => "11110100000000100000010000001111",
6385 => "11010110111101011111101011110101",
6386 => "11101111000000010000100111111101",
6387 => "11111010000000100000000111111010",
6388 => "11110100111101001111000000000001",
6389 => "00000100111100100000100111111110",
6390 => "11111110111100111111111100000010",
6391 => "11110111111101111111101111101110",
6392 => "11101011000000001110110000001011",
6393 => "11000111111101011110000111110110",
6394 => "11111010111100101111111100000100",
6395 => "11111011111110111111111011111100",
6396 => "00000110111111101111111011111101",
6397 => "00000010111111010000001000000001",
6398 => "00000101111111011111101000001010",
6399 => "11100111000001001111111011110101",
6400 => "00000101000000001110001111100100",
6401 => "11101110111111001111110000000000",
6402 => "00000011111110011111111100000010",
6403 => "11111101111111000000011000000000",
6404 => "00000110000000010000101111111111",
6405 => "11111100000000100000010000000000",
6406 => "00000111000000101111100000001001",
6407 => "11100100000000111111111011111010",
6408 => "00000011000010111100100011100111",
6409 => "11011110000001110000010100000101",
6410 => "00000101111111011110110111111001",
6411 => "00000011000000000000100111110111",
6412 => "00000011000001110000100011111010",
6413 => "00000011000001101111100100000000",
6414 => "00000001000001011111011100000100",
6415 => "11100101000011100000001111110111",
6416 => "11111101000001001110011011101010",
6417 => "11111001111111000000001000000001",
6418 => "11111100111110101110100111111100",
6419 => "00000100000000100000010111111010",
6420 => "00000110000001110000001011110101",
6421 => "00000100000001101111110111110000",
6422 => "00000001000011000000001100000010",
6423 => "11111111000101001111110100001011",
6424 => "11111000000001011111010111100000",
6425 => "00000000111101111111111100001010",
6426 => "00000101111101011101101011111101",
6427 => "00000100111111100000000111111111",
6428 => "00000101111110111111001111110101",
6429 => "00000100000000010000001011101111",
6430 => "11110100000000000000111111110101",
6431 => "11110101000001101111110000010011",
6432 => "11110101111110001111010011011101",
6433 => "11110111111110000000001100010100",
6434 => "11110011111110001101110111111111",
6435 => "11111100111110001111100000001000",
6436 => "11111001111111011111100111110110",
6437 => "11110111111111101111101011111010",
6438 => "11111110111111110000001011111000",
6439 => "11101100111100001111101000000100",
6440 => "11111111111110101111111011110111",
6441 => "11111110111111000000000100000101",
6442 => "00001010111111001110110011111010",
6443 => "11111110111101111111110000000001",
6444 => "11110110111111011111001011111011",
6445 => "11111110111010011111111111101110",
6446 => "11100001111101010000011111101100",
6447 => "11111011111001111111001000000111",
6448 => "11110110111111111111111000000010",
6449 => "11111101111011111111011111111111",
6450 => "11110101111110001111110000000011",
6451 => "11110001111011011111000111111011",
6452 => "11100101111010001110101011110010",
6453 => "11101101111010001111010111110011",
6454 => "11101010111000111111001111111111",
6455 => "11110111111001001110111111110101",
6456 => "11101001111001011111000100000011",
6457 => "11100100111110101101101011101110",
6458 => "11100000111001101110011111111001",
6459 => "11101001111101011111000011101010",
6460 => "00000001111111101111111011110101",
6461 => "00000001111101011111110111111010",
6462 => "11110010111110000000010011111100",
6463 => "11111101111111001111110111111101",
6464 => "11111110111101101111111111110111",
6465 => "00000011111100011111110111111110",
6466 => "11111111111101111111011011110111",
6467 => "11111001111101111111111111111101",
6468 => "11111000111111111111100011111110",
6469 => "11111001111100001111111011110110",
6470 => "11101011111010111111101011110000",
6471 => "11111011111100011111110111111000",
6472 => "11110001111100011111110111111011",
6473 => "11110101111110001111010011111011",
6474 => "11110011111111000000000111111000",
6475 => "11110011111110111111101011111100",
6476 => "11110011111010101110111111111010",
6477 => "00000001111001010000110111111001",
6478 => "11111000111111000000001111111110",
6479 => "11111001111100111111100011111010",
6480 => "11101000000001011111100000000011",
6481 => "11010101111100011101110111111000",
6482 => "11110010111101011110111111111101",
6483 => "11110100111101101111101011110011",
6484 => "11110010000110111111101111111101",
6485 => "11111011111000100000011011111010",
6486 => "00000010111110111111010100000100",
6487 => "11110100111011011111000111110010",
6488 => "11111011000110001110110100010001",
6489 => "10110111111110011111101011111000",
6490 => "00000000111100010000001011111011",
6491 => "11110000111101111111110111111010",
6492 => "11110100000011001110111000000101",
6493 => "11110010111100100000001100000010",
6494 => "00000100111110101110100100000100",
6495 => "11101000111100111111100111100100",
6496 => "11111101000000001100100000000011",
6497 => "10101100111111111110010011101010",
6498 => "00000001111101010000010000000010",
6499 => "11110011111110001111110011101001",
6500 => "11111100000110011111010111111100",
6501 => "11111000111000010000111111111000",
6502 => "00001111111111001110101000001001",
6503 => "11110000111101001111010011110001",
6504 => "00000001000011011100110011110000",
6505 => "11110100000001011110010111101110",
6506 => "00001011111010001111000100000011",
6507 => "11110011111111011111111111100101",
6508 => "11110111000011101111111111110101",
6509 => "11111010111001000000010011111110",
6510 => "00010001111110001111000100010000",
6511 => "11101111111010101110111100000011",
6512 => "00000110000110011100010011110011",
6513 => "11101110000001101111110000000000",
6514 => "00001010111110001110001000000111",
6515 => "11101110111111001111111011111100",
6516 => "11111111000001111111111011110101",
6517 => "11111101111101111111001111111010",
6518 => "00010100111111111111111100001011",
6519 => "11111000000001011111101000011111",
6520 => "00000000111111111100000111011010",
6521 => "11111000000001010000000000010100",
6522 => "11111110111101101011011111111010",
6523 => "11111010111111011111010100000101",
6524 => "00000000000100111111110111100001",
6525 => "11110100000010101110100111110101",
6526 => "00001111111110010000010000010111",
6527 => "00001001111101101111100000100101",
6528 => "11111111000000101110001011011110",
6529 => "00010001000001010000111000001101",
6530 => "00000001111110111100010011111000",
6531 => "11110111111110111111010000000011",
6532 => "00000101111111000000100111110111",
6533 => "11111000000100011111001111111001",
6534 => "00010010111111100000010100001111",
6535 => "00000011111111111111110000101011",
6536 => "11111111111100100000100011010101",
6537 => "00001001000001000001000100001110",
6538 => "11111011000010101111010111111010",
6539 => "11111001000001101111101000001101",
6540 => "11110111111111001111011111111110",
6541 => "00000100000001110000000111111001",
6542 => "00000010000100100000100000000000",
6543 => "11110111000000110000000100010001",
6544 => "00001001111111010000000100000000",
6545 => "00000111000001010000111000010011",
6546 => "00000110000010001111110111111010",
6547 => "00000000111111001111111000001010",
6548 => "11111101000000011111010011111111",
6549 => "00000011000001110000000011101111",
6550 => "11101101000010101111101111111010",
6551 => "11111110000011011111011111110100",
6552 => "11111100000000000000110011100101",
6553 => "00010000111111110000001111110010",
6554 => "11111100111110000000110011111000",
6555 => "11111101111101101111010100000001",
6556 => "11101001111100011111001111111111",
6557 => "11101111111100101111001111111010",
6558 => "11101010111111111110011111111101",
6559 => "11111000111100001111100111111111",
6560 => "11110001111010100000100011101001",
6561 => "11110101000000111110100011100110",
6562 => "11101011111010110000001111111011",
6563 => "11110001111111101111011011101011",
6564 => "11111101000000001111101011111110",
6565 => "11110111000000001111101111110110",
6566 => "11100100111110001111011011110111",
6567 => "11111011111111101111100011111011",
6568 => "00000011111110110000001011111101",
6569 => "11111111111101011111111011111011",
6570 => "00000100111111100000001011111100",
6571 => "00000001111110101111101011110111",
6572 => "11110111111110111111011111111001",
6573 => "11011010111101101111010111101000",
6574 => "11101111111101101101001111111000",
6575 => "11111010111101101110111111100111",
6576 => "11101101111000000001000100000101",
6577 => "00010010110110010000011111010101",
6578 => "11101100111110011110111011110111",
6579 => "11110011111110001111000011000010",
6580 => "11110100110110111111110100001001",
6581 => "11100111111001011110100111111111",
6582 => "11110100111110001110100111111100",
6583 => "11111000111011011111010111101101",
6584 => "11101010111101000000000100000001",
6585 => "00001000111111011110111011110001",
6586 => "11101101111111000000101011111011",
6587 => "11111001000000001111110011101101",
6588 => "11101010000101101111011011111100",
6589 => "11110010111100101111101111111010",
6590 => "00001010000001101111001100000011",
6591 => "11111001000001011111010111110110",
6592 => "11110111000010101111011011110101",
6593 => "11111100000001011111010011110010",
6594 => "00001001111101001110101100000000",
6595 => "11101111111111111111110011101100",
6596 => "11110101000011101111000011111010",
6597 => "11100000111001101111010111111110",
6598 => "00001010111111101110101000001100",
6599 => "11110101111101011111100111110100",
6600 => "00000100000100101100111111111001",
6601 => "11101011000001000000001011101010",
6602 => "00001011111011111110100111110111",
6603 => "11110001111110100000001111100011",
6604 => "11110100000111101110101011110011",
6605 => "11101101111000001111010111101111",
6606 => "00010001111111011110110000001010",
6607 => "00000000111001101111010100000011",
6608 => "11111100000100011101001011111111",
6609 => "00010011000010101111100111110000",
6610 => "00000000111111001101111011111001",
6611 => "11110010111111011111010011110001",
6612 => "11101011000101011111001011111001",
6613 => "11110000111011111111001011111000",
6614 => "00001100111110001110110000001111",
6615 => "00000101111100001111100100000110",
6616 => "00000010000000101101101011101111",
6617 => "00011010000000010000010011110101",
6618 => "00001101111101101110001000001010",
6619 => "11110101111111001111011111101101",
6620 => "11111011000110001111100011110001",
6621 => "11110010111100111111000111110111",
6622 => "00010000111111001110101000010000",
6623 => "00010001111100011111010100001000",
6624 => "00000001111111101110110111100010",
6625 => "00011111000001110000010011110100",
6626 => "11111111111111001100111111111100",
6627 => "11110100000000001111010011101101",
6628 => "11111010000010001111101111111001",
6629 => "11110100000001101111011100000001",
6630 => "00001101111110111111001100001110",
6631 => "00010010111110001111100100001010",
6632 => "11111111111111100000000011110011",
6633 => "00000100000000100000011011110100",
6634 => "11111001000001011111111100000101",
6635 => "11111111000000011111101011110110",
6636 => "11111010000001111111011111111110",
6637 => "00000100000000010000001000000011",
6638 => "00001010000000010000011000001001",
6639 => "11111111111111001111100100010110",
6640 => "00000010000000011110111011110000",
6641 => "11111110000011010000001000000101",
6642 => "00000011111111111111000111111001",
6643 => "00000000111110011111101100001000",
6644 => "00000001111111101111111100000111",
6645 => "00000100000001000000100111111101",
6646 => "00000101000000000000111100001000",
6647 => "11111010000000001111101100001010",
6648 => "00000111111111011111110000001101",
6649 => "11111101000001000000100100001010",
6650 => "00000101111111111111001011111100",
6651 => "00000001111110111111111100000110",
6652 => "11111110000000100000010011111101",
6653 => "00000000111011100000010111111100",
6654 => "11110100000000100000100111111011",
6655 => "11111101111001101111011111111101",
6656 => "00000001000001110000010000010111",
6657 => "00000011000000000000000100000101",
6658 => "11111111000010000000001111111101",
6659 => "11111110000001010000000011111111",
6660 => "11111101111100100000000111111101",
6661 => "11111011111111101111101111111110",
6662 => "11101010000001011111011000000001",
6663 => "11111110111110100000001011111010",
6664 => "00000000111101001111110000000001",
6665 => "11110101111111001111011011111000",
6666 => "11111101111110100000010011111100",
6667 => "00000001000010010000000011110100",
6668 => "11111101111111001111111100000000",
6669 => "00000001111111110000001000000010",
6670 => "11101010000000000000001011111011",
6671 => "11111001000000100000001011111110",
6672 => "11111101111101110000010111110111",
6673 => "00000101111111111111111011111111",
6674 => "11111111000000110000000011111100",
6675 => "00000011111111010000000111111111",
6676 => "11111111111111000000000100000111",
6677 => "00001110000010011111011100000101",
6678 => "00001010000001000000010100001101",
6679 => "11111010000001101111101100001000",
6680 => "00000001111111010000010000001010",
6681 => "00000100000001110000101000001101",
6682 => "11111110000010100000100111110110",
6683 => "00000111000010110000010100001101",
6684 => "11111010000011111111101000000101",
6685 => "11111111000001000000010000000110",
6686 => "11100100000000100000001111111011",
6687 => "11111010000010110000001111111011",
6688 => "00000110000011000000111011101101",
6689 => "00010001111010000000001011111010",
6690 => "00001011111101010000100111111100",
6691 => "00000000111110010000001111111000",
6692 => "11101110000101001111100111101101",
6693 => "11110000111001101111010011101110",
6694 => "11110110111010001111011111111101",
6695 => "00000010111100111110110111111011",
6696 => "11101111000011110000000111111101",
6697 => "00001000000000101110100111111100",
6698 => "00000100111110101111111000000001",
6699 => "11100110111010011110111011110000",
6700 => "00000010000000011111101011100110",
6701 => "11111100000000110000001000000001",
6702 => "11110111000000101111101000001011",
6703 => "00001001000000111111010000001000",
6704 => "00000010000001111111110000001010",
6705 => "11110010000001010000100011111100",
6706 => "00001000111111111101110000000001",
6707 => "11111100111110001111011011111011",
6708 => "11110100000011001110110011101100",
6709 => "11110111000000101111101011101111",
6710 => "11110010111100001111101011111101",
6711 => "00000101000000001111101011111100",
6712 => "11110101000001101111101100010000",
6713 => "11111111111100001110111011101110",
6714 => "11111000111011101100100100000000",
6715 => "11110110111011111111010011110100",
6716 => "11111110111101111111101011101001",
6717 => "11110001111101001111011111110101",
6718 => "11111110111010111111100000000011",
6719 => "00000111111100101111001100000101",
6720 => "11111010111110001111101011111100",
6721 => "11101001000000010000001011111010",
6722 => "00000001111101111101100000000011",
6723 => "11110000111111001110110111111001",
6724 => "11110000111111101111000111101001",
6725 => "11110101111100101111100111110010",
6726 => "11110100111010001111110000000001",
6727 => "00001010111100011111100000000111",
6728 => "00000010000000101111111000001101",
6729 => "00000001111100101111110011111010",
6730 => "11110110111011001110110000000010",
6731 => "11101100111110001111000011110100",
6732 => "11111000111101001111110011110000",
6733 => "11111001111011111111110111111101",
6734 => "11010110111010111111110111101100",
6735 => "00001011111110001110110100001000",
6736 => "11111000111111000000101100000100",
6737 => "11101001111000111111001011111010",
6738 => "11111000111010110000000000000101",
6739 => "11101010111010111111111011110110",
6740 => "11110110111011111111101111110111",
6741 => "11110011111010111111100011110011",
6742 => "11100111111010110000000111110000",
6743 => "11111101111010001111010111111100",
6744 => "11101101111111111110101100011100",
6745 => "11011110111100111111010111110111",
6746 => "11101101000001011110011111111111",
6747 => "11101111111101011111010011110001",
6748 => "11111111111000011111111111111010",
6749 => "11110111111101101111100111111100",
6750 => "11110001111101110000000111110101",
6751 => "11111001111010001111100000000011",
6752 => "11111010111010101111100011111110",
6753 => "11010000111100010000011100000010",
6754 => "11110110000000111111001011111111",
6755 => "11110010111101111111111000000001",
6756 => "11110000111111101111010000000010",
6757 => "00000001111011110000000100000000",
6758 => "11101011000000111111101100000011",
6759 => "11110111111100011111110111110111",
6760 => "11110000111111010000011100000100",
6761 => "11111000000000111111011011110100",
6762 => "11110011111101011111101111110111",
6763 => "11111000111110101111110111110101",
6764 => "11111110111100110000000111111110",
6765 => "11111011111111101111110100000001",
6766 => "11101010000000011111101111111100",
6767 => "11111000111110010000001011111001",
6768 => "11111110111100100000010011111100",
6769 => "11111110000000101111110111111001",
6770 => "00000001111110110000001011111100",
6771 => "00000101000001000000011011111101",
6772 => "00000000000000000000000000000000",
6773 => "00000000000000000000000000000000",
6774 => "00000000000000000000000000000000",
6775 => "11111100111111100000001100000011",
6776 => "00000010111111001111110100000010",
6777 => "00010010000000011111100100000010",
6778 => "00000100111111001111110111111100",
6779 => "00000001000001011111110111111110",
6780 => "11111001000000000000000100000001",
6781 => "00000001111111000000001100000000",
6782 => "11111101111111011111110100000100",
6783 => "11111001000011111111111000000000",
6784 => "00000011111111111111011011111101",
6785 => "00010011111111100000000000001011",
6786 => "00000001111111111111101111111010",
6787 => "00000100000001100000010000000111",
6788 => "00001010000000001111100100000001",
6789 => "00000000111111100000111100000001",
6790 => "11111010000000011111111100000011",
6791 => "11111010000100011111101011110000",
6792 => "00000000111110001111011111110101",
6793 => "11110001111100111111110011111011",
6794 => "00000100111100111111101111111100",
6795 => "11111000000011110000100111111111",
6796 => "00001010111100001111000011111110",
6797 => "11111110111110000000110000000100",
6798 => "11111000111101001111110111111111",
6799 => "11101110111110000000000111110101",
6800 => "00000011111100111111101111111011",
6801 => "00000000111110001111101000000010",
6802 => "00000001111100101111101100000000",
6803 => "11101111000001110000001000000011",
6804 => "11110110111100111111110100000001",
6805 => "11110100111111101111010000000100",
6806 => "11110110111101111111101011111110",
6807 => "11101100000000000000001100000000",
6808 => "00000000111011001111110011111010",
6809 => "11111101111100111111110000000000",
6810 => "00000000111010101111011111111010",
6811 => "00000110111011110000100100000001",
6812 => "00000001111011001111110111111000",
6813 => "00000010111111000000000000000100",
6814 => "11110010111111001111111111111011",
6815 => "11110111000001011111001111110100",
6816 => "11111111111000011111101111110100",
6817 => "11110101111100001111100011111101",
6818 => "00000101111010111110110111111101",
6819 => "11110110000010000000000011110111",
6820 => "11111100111000001111011111111100",
6821 => "11111110111101001111110111111111",
6822 => "11110100111100001111001111111110",
6823 => "11101010000000011110110011110100",
6824 => "11111010111000111111110111110101",
6825 => "00000101111101001111011000000100",
6826 => "00000111111011001111101111111100",
6827 => "11110111111101011111111000001000",
6828 => "11111101111100111111100011110010",
6829 => "11111011111110111111100000000101",
6830 => "11111011111110001111100011110111",
6831 => "00000110000000101111001011111000",
6832 => "11111111000001001111011011111110",
6833 => "00001001111110001111011000000111",
6834 => "00000100000011000000000111111101",
6835 => "11111000000001110000001100000111",
6836 => "11111010000100001111110111111110",
6837 => "11111000111111011111100100000100",
6838 => "11111101111111001110111011111000",
6839 => "00000000000000100001000000001010",
6840 => "11110010000001101111101000000010",
6841 => "00000101000001101111010000010111",
6842 => "11111100111111111111110111111110",
6843 => "00010001111001000000011100010010",
6844 => "00000100000001000000111111110110",
6845 => "00000010000011111111111000000000",
6846 => "00001000000100001111110111111001",
6847 => "00000111000101000001000100000100",
6848 => "11111101111110001111011011111100",
6849 => "11110110111111001111011111111111",
6850 => "00000111111111011111110011111110",
6851 => "00000011000101010000110100000100",
6852 => "00001111111110001111011111111001",
6853 => "00001001000000000000110000000101",
6854 => "11111001000000100000000100000100",
6855 => "11111010000001101111101011111111",
6856 => "00000100111110011111111000000001",
6857 => "11111010111100110000000000000010",
6858 => "00000110111111011111101111111101",
6859 => "00000001111111000000010011111101",
6860 => "00000100111110010000101011111101",
6861 => "00001011000001010000011100000101",
6862 => "11110111111111110000100111111111",
6863 => "11111110111110011111111011111010",
6864 => "00000110111111001111110111111001",
6865 => "11110010111101111111101111111001",
6866 => "11111101111111011111011011111010",
6867 => "11111101111110011111000111101111",
6868 => "11101100111101111111001111111101",
6869 => "11110010111110101110111100000110",
6870 => "11111011111111011111011111111111",
6871 => "11111111111111011111110111111111",
6872 => "00000000111111111111101011111111",
6873 => "00000100000001011111111000000111",
6874 => "00000011111111011111111011111101",
6875 => "00000101111111011111101000000000",
6876 => "11111010111111001111111100000101",
6877 => "11111011000000111111100000000011",
6878 => "00000000111111001111100111111111",
6879 => "11111101000000101111101100000000",
6880 => "00000001111111111111100011111111",
6881 => "00010010111111111111101000001110",
6882 => "00000010111111101111101011111011",
6883 => "11111100000010001111110000001001",
6884 => "11110011111101101111101100000010",
6885 => "00000010111111101111110000000001",
6886 => "11111011000000101111111011111111",
6887 => "11110001000100001111101011101011",
6888 => "00010010111010110000001011111000",
6889 => "11111000111110011111100011111110",
6890 => "00000110111101011111001011111111",
6891 => "11110111000011011111101111110111",
6892 => "11110100111011001111010011111000",
6893 => "11111100111011001111110000000011",
6894 => "11110111111011001111101000001010",
6895 => "11101110000010001111011011110110",
6896 => "00000000111101100000011111111011",
6897 => "11110000111110010000011011110011",
6898 => "00000000111011001111100011110110",
6899 => "11101001000100111111001011110001",
6900 => "11101101111100011111100011101111",
6901 => "11110011111110111110110100000011",
6902 => "11110100111101101111010011110110",
6903 => "00001000111001101110110011111000",
6904 => "11100010111001101111100111111001",
6905 => "00001101111011101111000100001100",
6906 => "11111110111111111111110011111111",
6907 => "11110001111100001111101000000101",
6908 => "11101101111101111111111000000000",
6909 => "11110111111111011110110000000101",
6910 => "11111010111111001111000011101010",
6911 => "11110111111001010000100100000111",
6912 => "11101000111101000000001100000011",
6913 => "00000001111110011101111100001001",
6914 => "11111101111110101111111011111000",
6915 => "00000111111100100000001100000111",
6916 => "00000011111111001111111111111011",
6917 => "11111001000001000000100000000010",
6918 => "11111101000011000000000011010010",
6919 => "11110100110110010000001011111110",
6920 => "11011011111010100000011011111100",
6921 => "11110110111100101100001011110101",
6922 => "11110001111010001111011111100010",
6923 => "11111010111001000000000111111100",
6924 => "11110110111101001111011011001001",
6925 => "11111010111101111111110000000101",
6926 => "11110100111110111111111011000011",
6927 => "11111110110100101111100011111000",
6928 => "11101000111011110000100100000110",
6929 => "00000000111101011110011100000010",
6930 => "11110111111001010000000111100111",
6931 => "00000010111101101111011111111010",
6932 => "11101111000000011111010111101011",
6933 => "11111101111111001111110011111110",
6934 => "11110101000001000000010011101101",
6935 => "11110100000000011111111011111100",
6936 => "11111100111101100000010100000100",
6937 => "00001101111111101110111100001100",
6938 => "00000001111100110000010011110011",
6939 => "00001000000101101111101000000111",
6940 => "11110010000010011111110111101000",
6941 => "00000100000001000000000011111100",
6942 => "00000010000001010000000011110111",
6943 => "11111010111111110000001100000100",
6944 => "00000100000000000001000100001000",
6945 => "00001000000001111111001100001110",
6946 => "00000001000000010000010111111010",
6947 => "00010001000010111111101000000000",
6948 => "00000001000011000000100111101001",
6949 => "00010001000001000000010100000110",
6950 => "00001011000001000001000011111110",
6951 => "11110011000011000000001111111010",
6952 => "00010101000000010010000100000001",
6953 => "11110111000010100000111011110010",
6954 => "00000010000001000000010011110100",
6955 => "11111001000110001111100111110001",
6956 => "00000011111110011110110000000101",
6957 => "00001101111101011111100000000010",
6958 => "00000100111101100000100000001101",
6959 => "11110001111111010000110011111010",
6960 => "00010000000001000001001000000100",
6961 => "00011011000001000000001000010111",
6962 => "11111011111111101111110111110110",
6963 => "11111110000100101111001000010011",
6964 => "11110001000010101111010011111111",
6965 => "00000010111111111111011100000001",
6966 => "00000001000010110000001011111110",
6967 => "11110011111111110000100100000000",
6968 => "00001001111111010000101100000000",
6969 => "00000001000011100000101100001011",
6970 => "00000001111111111111100011111001",
6971 => "11111100000000101111100100011001",
6972 => "11111011111111101111010100001001",
6973 => "00000001111101001111100000000100",
6974 => "11111111000001110000101000001100",
6975 => "00000010000010110000011000001000",
6976 => "11111111111110011111110000000110",
6977 => "00001110000010101111101000001101",
6978 => "00000101111111111111111100000001",
6979 => "00000000000001110000011000001100",
6980 => "00000101111111010000001011111111",
6981 => "00000110000000100000011000000110",
6982 => "00000101000001100000100000000001",
6983 => "11101000000001001111100011101111",
6984 => "00001000111010011111101111110001",
6985 => "11111111111110000000110100000110",
6986 => "00000001111010011111001000000110",
6987 => "11111111000001100000000100000000",
6988 => "00000110111110001110000100000100",
6989 => "00001001111011100001001000000110",
6990 => "11110010111011101111110000000111",
6991 => "00000110000100011111000111110011",
6992 => "11101011111110110000001011110011",
6993 => "00000101111111101110110100000000",
6994 => "00000100111110011111100111110011",
6995 => "11110101000100101111001011111110",
6996 => "11110001111111001111000111110011",
6997 => "11110111111101011110001100000011",
6998 => "11111010111111011111010111100101",
6999 => "11111000000010001111110111111110",
7000 => "11001100111110001110000011111011",
7001 => "11111000111100101101011111111001",
7002 => "11111111111101111111110011110000",
7003 => "11111100111001001111100111111101",
7004 => "00000010111101001111110011101000",
7005 => "11111110111110111111100100000001",
7006 => "11111101111111101111011111010111",
7007 => "11110111000000000000001000000011",
7008 => "11011000111111111101001100000110",
7009 => "11111010111111011100100100001000",
7010 => "11111000111100101111110111111001",
7011 => "00000010111100101111111100000000",
7012 => "11110110111111000000010111110000",
7013 => "00000010000000011111101111111101",
7014 => "11111000000000101111111111001111",
7015 => "11111001111110000000001000000100",
7016 => "11101110111110111110110011111001",
7017 => "11111110111111111110000000000110",
7018 => "11110010111111100000000111111101",
7019 => "00000111111100010000000111110000",
7020 => "00000000000001001111101000000100",
7021 => "00001000111110001111011100001010",
7022 => "11111111111111101111110111110100",
7023 => "11101110111011101111011100001000",
7024 => "11111010111101100000111011111100",
7025 => "00001001111111111110010100000010",
7026 => "11100000111110101111111111110011",
7027 => "00000100000101001111100011110011",
7028 => "11110111000010101110110011111001",
7029 => "00000100111100111111111000001100",
7030 => "00001000000000011111110011110010",
7031 => "11101011111001001111111100000101",
7032 => "11111111111101000001100100000110",
7033 => "00000100000001001111101011111010",
7034 => "11100100111101011111100011101101",
7035 => "00000010000000011111010011111010",
7036 => "11111011000000011111000111101111",
7037 => "00001110111100101111101100001001",
7038 => "00000000111111100000000100000011",
7039 => "11101101111011011111011000000110",
7040 => "00001010111100010001101000000011",
7041 => "00001010000001000000000000000000",
7042 => "11100011000000001111110011111000",
7043 => "00000100000011001111100000010001",
7044 => "11110101000010101110011000000001",
7045 => "00000101111101111111101100000011",
7046 => "00000001111111101111111100000001",
7047 => "11111111111111100000000100000100",
7048 => "00001001111101000010000000000110",
7049 => "00000110000001011111111011111111",
7050 => "11110010111110110000000011101001",
7051 => "11111011000101111111110000011111",
7052 => "11111001000001111111010111101110",
7053 => "00001100000000000000010100000111",
7054 => "00000111111101100000001011111110",
7055 => "11101111000000011111110100001011",
7056 => "00010000111010010010111000000101",
7057 => "00010110111111000000111111111111",
7058 => "11110000111011111111101011101001",
7059 => "11111111000101101111111000110110",
7060 => "11110001111111011110100011111010",
7061 => "11111110000000011111110100001010",
7062 => "00000001111111011111111100001010",
7063 => "11101110111100111111010000001110",
7064 => "00010011110111010010111000000100",
7065 => "00100111111101100001100100100010",
7066 => "11111111111101001111000011110010",
7067 => "11100100000101011111111101000011",
7068 => "11110111000010101110001000000010",
7069 => "11101100111110010000100000001011",
7070 => "11110100000000001111001100001010",
7071 => "11111001111100100000010100001111",
7072 => "00010111111101000001010000001000",
7073 => "00000101000010010001101100000101",
7074 => "11110111111110011111100100001001",
7075 => "11111100000000001111010000101100",
7076 => "11101111000010001111011000010110",
7077 => "00000001111101101111111000000110",
7078 => "00000100000000001111111000010111",
7079 => "11111111000000100000101000001111",
7080 => "00001110111110110000011100001010",
7081 => "00010111000101111111111000010001",
7082 => "11111110000011100000101111110110",
7083 => "11111111000010011111101100010100",
7084 => "00000000000010011111101111111011",
7085 => "00000110111111011111101100000100",
7086 => "00001001000010000000100100000001",
7087 => "11101011000000111111001011100011",
7088 => "11101110111001010000000111101011",
7089 => "11011101111011011110011111101110",
7090 => "00000101111001011111000111110011",
7091 => "11111001000011001111100111110001",
7092 => "11101110110111101110111011101000",
7093 => "00001001111001101111000000000110",
7094 => "11101110111001011111010111100110",
7095 => "11101101111111101111001011111001",
7096 => "11101101111001111111000011110011",
7097 => "00001000111011011111001100000011",
7098 => "11111111111011011111010111111111",
7099 => "11111011111110111111000000000010",
7100 => "11100100111111111111000011111110",
7101 => "11111001111111001111001000000101",
7102 => "11110000111111001111101111110110",
7103 => "00000111000011110000010011110110",
7104 => "11010111000000011101001000000010",
7105 => "00000011000000101101110100000100",
7106 => "11110101000010001111110111111111",
7107 => "00000101000000011111000111101110",
7108 => "11110111111110100000101111111100",
7109 => "11111111111111101110111000000000",
7110 => "11111101000001001111101111100000",
7111 => "00000001000010110000110111111100",
7112 => "11010100000010001100110000000001",
7113 => "11111010000000011101001011111110",
7114 => "11110100000010110000011011110110",
7115 => "00001011111011111111010011100001",
7116 => "00000010000000100000101011111010",
7117 => "00000110111110111110100000000100",
7118 => "00000101111111110000010011100011",
7119 => "11111011000101011111101111111110",
7120 => "11101101111100001110000011111100",
7121 => "00000000111111001110001011111010",
7122 => "00000110111111000000000111111110",
7123 => "00000111111111001111110011011110",
7124 => "00010010000000011111011000000111",
7125 => "00000001111101111111000100001110",
7126 => "11111101111111101111101011110001",
7127 => "11111101000100000000100111111111",
7128 => "11111011000001001111011111111111",
7129 => "00000100000001111111000100000101",
7130 => "11110010111111010000001100000100",
7131 => "00001110111111111111011011100000",
7132 => "00001101000001010000101100001001",
7133 => "00001011111110011110111100010000",
7134 => "00000010111111100000011000000001",
7135 => "11111100111111110000000011110111",
7136 => "00000001111101000000100100000100",
7137 => "11110111111110111111111111101001",
7138 => "00000011111101100000011000001011",
7139 => "00000100000000011111000111101000",
7140 => "11111101111111101110110000000011",
7141 => "00000011111101001110110100101001",
7142 => "00000010111101001111111100000011",
7143 => "11111011110010001111111000000111",
7144 => "00001110000000000001101000000011",
7145 => "11100101000000010000111111001111",
7146 => "11111001111111000000010000011000",
7147 => "11111111111011110000110111111011",
7148 => "11110111111111101111000100001110",
7149 => "11101010111111011111100100101000",
7150 => "00000011111101001111110000010010",
7151 => "11110110110100001111101000001000",
7152 => "00010101111101000010000111111110",
7153 => "11001101000001000001010110110101",
7154 => "11101111000010001111101111111011",
7155 => "00000000000000010001100000011111",
7156 => "11111001111101101110011100000110",
7157 => "11111101111100000000000000011001",
7158 => "00000011111010001111001000010000",
7159 => "11111100110101011111010000001101",
7160 => "00100010111001100011001100000010",
7161 => "11101011000010000010101111001000",
7162 => "11100111000001011111110011111101",
7163 => "11111100000011000010000000111001",
7164 => "11111110111110001101111100010011",
7165 => "11110101111011100001001000010001",
7166 => "00000100111010001111111000011101",
7167 => "11111000110101011111101100001100",
7168 => "00011111111001100011000100000100",
7169 => "11101110000001010001101011011111",
7170 => "11110000000001111111110111101011",
7171 => "11101000000001010001011100111100",
7172 => "11110110111110001101101100001010",
7173 => "11100111111011000001010100001100",
7174 => "11111011111011111110111100011001",
7175 => "11111100111001010000011100011000",
7176 => "00001001111101000000111000000010",
7177 => "11111010000010010000110111110010",
7178 => "00000000000000111111100111110010",
7179 => "11111110111101100000101100101110",
7180 => "11110010000001011110111000000110",
7181 => "00000100111111000000111111111111",
7182 => "00000011000000010000001000000110",
7183 => "00001101000010000000111000011011",
7184 => "00010011000000110000100000001110",
7185 => "00010110000010100000110100000101",
7186 => "00000111000011100001000011111000",
7187 => "00000001000010010000110000101000",
7188 => "00000110000010110000011000010100",
7189 => "00000110000101110001100100000011",
7190 => "00001110000100000001001000001001",
7191 => "11101100111111101111010011101010",
7192 => "11100001111001101111010011101100",
7193 => "11011001111010101101101011101100",
7194 => "00000001111010111110110111110010",
7195 => "11110010000010001111110011110110",
7196 => "11101011111000001110110111100110",
7197 => "11110110111011101110100100000101",
7198 => "11110001111010111110101111011100",
7199 => "11111000111101000000000100000000",
7200 => "11110000111111011101101111110111",
7201 => "00000001111111011110110000000011",
7202 => "11111101111110111111010100000110",
7203 => "00000000111000001111111000000111",
7204 => "11011111111111110000010011110101",
7205 => "00001001000000110000011000000001",
7206 => "11110111111111001111111111110011",
7207 => "00001001000110010000000011111111",
7208 => "11100010000011001101101011111111",
7209 => "00000010000000011110111011111110",
7210 => "00000001000001010000010111110001",
7211 => "00000000111110011110111111100100",
7212 => "11111001000001010000011111110100",
7213 => "00000000000010001111100011111011",
7214 => "00000011000000100000011111101010",
7215 => "00001100000101010000011011111101",
7216 => "11101111000110101101010100000011",
7217 => "00001001111111001111001100000010",
7218 => "00001000000000100000010111111101",
7219 => "00000010111010111110001111011100",
7220 => "00000010000010010000100000000011",
7221 => "00000100000010111110011100000010",
7222 => "00000100000001010000011111110111",
7223 => "00000010000100111111111100000010",
7224 => "11110010000010101101100100000110",
7225 => "00000000000010101110111000000100",
7226 => "11110000000010110000010100000100",
7227 => "00001100111110111111100111100010",
7228 => "00011101000000110000100000000010",
7229 => "00010001000001111111010100000110",
7230 => "00000100000001010000011011110111",
7231 => "00001000000011100000111000000101",
7232 => "11111010111111111111110000000010",
7233 => "00000010000001001111101000000101",
7234 => "00010100111111000000011000001101",
7235 => "00001010111110100000010011011010",
7236 => "00100000000010110001010000000111",
7237 => "00000011000010001111101000001010",
7238 => "00000010000010000000000111111101",
7239 => "00000100111111100000101111110110",
7240 => "00000010111100111111111011111100",
7241 => "11110011000001100000000111100101",
7242 => "00011111000000100000000000011010",
7243 => "11111111111111110000001011101011",
7244 => "00011000111111101111010000000110",
7245 => "11111111111111101110111000100100",
7246 => "00000110111111011111111000000100",
7247 => "11110011110010110000011111111011",
7248 => "00000011111101010000101011111010",
7249 => "11000110000000110000111110110111",
7250 => "00011100111111111111010100101001",
7251 => "11111111110111000001100011011011",
7252 => "00001110111001101110110000010000",
7253 => "11110001111010011110111100110000",
7254 => "11111111111101001111001000001010",
7255 => "11111010110010111111100011110011",
7256 => "00010011111110010000111011110000",
7257 => "10100110000001000010010110011000",
7258 => "00010111000000101111011100110001",
7259 => "11110111110101010010001011011001",
7260 => "00011100111010101111000100100011",
7261 => "11101110111011011111001000011110",
7262 => "00000011111011001111010100100011",
7263 => "11110001110001011110110111111100",
7264 => "00010100111110010010000011101000",
7265 => "10111101000001010010000010010110",
7266 => "00010010000010111111100100001110",
7267 => "11100011111010010010010011101111",
7268 => "00011001111010111101101100011010",
7269 => "11101001110111101111111100011000",
7270 => "00000000110101001110111100011110",
7271 => "11111011101101011110110000001011",
7272 => "00001101111111100001011011110001",
7273 => "10111100111101010001010111000000",
7274 => "00000101000000101111110100000100",
7275 => "11100101110111110010001011111010",
7276 => "11111111111011011110010000001101",
7277 => "11100011111001000000000100010000",
7278 => "11111100111010001111000000010101",
7279 => "00000000110111000000010000010010",
7280 => "00010101111111000000110100000111",
7281 => "11011011000100000001100111010100",
7282 => "11111101000001110000101111111011",
7283 => "11111001111100110000111100010011",
7284 => "11110101111101101111110000010011",
7285 => "11111100000011100000100100001001",
7286 => "00010100111110010000101000010100",
7287 => "00010000000011100000110100010011",
7288 => "00011001000110010001101100010011",
7289 => "11111110000110100001011111111000",
7290 => "00000010001000110000110111110010",
7291 => "00001001000011110001011000000101",
7292 => "00010110000010010000110100001101",
7293 => "00001110000011100001010011111111",
7294 => "00010101000100110000100000010110",
7295 => "11110100000001011111110011110100",
7296 => "11100111111100101111011011110111",
7297 => "11110000111110001110000111111011",
7298 => "00000011111100001111010011110100",
7299 => "11111010000001101111100100000011",
7300 => "11110110111100011110101111101100",
7301 => "11111010111101001110111000000010",
7302 => "11110101111101001111010111100001",
7303 => "00001010111100110000000111101101",
7304 => "11101100000000111110111111111100",
7305 => "11111000111110101111110011111001",
7306 => "00001011000001101111110011111111",
7307 => "11111000111010111110010111101110",
7308 => "11010110111111011111110011111111",
7309 => "11110111111110001110010000000001",
7310 => "11111001111110101111110011111001",
7311 => "00001110000001000000100011110110",
7312 => "11101010000011001110010100000011",
7313 => "11111110111110011111011111111100",
7314 => "00000110000010000000001100000101",
7315 => "00000000111010011101110011100100",
7316 => "11111001000000010000100100000101",
7317 => "11111110000000101110000000000100",
7318 => "00000000111110010000010011111111",
7319 => "00000100000001110000010111111100",
7320 => "11101111000010111110010111111101",
7321 => "11111001000000011111011011111100",
7322 => "00010110111111101111111100001000",
7323 => "00000101110111011110001111100001",
7324 => "00010110000000100000001000000010",
7325 => "00000001000010001111001000001010",
7326 => "00000000111111100000100111111111",
7327 => "00000000000101000000010000000001",
7328 => "11110111111101110000000000000100",
7329 => "00000111000000111111110100001000",
7330 => "00001100111111100000010100000100",
7331 => "00001000111110001110010111101010",
7332 => "00010100111111110000010000000110",
7333 => "00001101000010011111100100001010",
7334 => "11111111000011100000111011111001",
7335 => "11111111000010010000100000000111",
7336 => "11110001111011111111100100000011",
7337 => "11111111111111111111010100000010",
7338 => "11111101111101110000100000000001",
7339 => "00001000000010101111011111100001",
7340 => "00001110000001111111010011110011",
7341 => "00000010000001001111000000010011",
7342 => "00000110000011010000010111110111",
7343 => "11111010000000001111111000000110",
7344 => "11111111111101111111110011110110",
7345 => "11111001111111101111111011100101",
7346 => "00001111111110001111110100010111",
7347 => "11111110111110110010000111101100",
7348 => "00011100111111011110101100000101",
7349 => "00000011111111100000011000010110",
7350 => "00000000111110011111110000000101",
7351 => "11111101110111010000000011110111",
7352 => "00001110111110100000110111101101",
7353 => "11000011111110110001001010110010",
7354 => "00100000000000011111010100100101",
7355 => "11111011111001110001100011011111",
7356 => "00010011111001011110110100001110",
7357 => "11111011111100111111111000011010",
7358 => "11111101111110111111100100001110",
7359 => "11111010110111000000010011110000",
7360 => "00000010000001011111101011101011",
7361 => "11000001111110010001011110110001",
7362 => "00100011111111001111110000101111",
7363 => "11111100101111110001011110111100",
7364 => "00011001111010011111011000011111",
7365 => "11110010111101001111100000100001",
7366 => "11111001111100011111001100010000",
7367 => "11101101111001011111010111101111",
7368 => "11111110111111011111110011100111",
7369 => "10110101111100110001011110100111",
7370 => "00100000111110111110100000100101",
7371 => "11110100110101000001101111011000",
7372 => "00011010111011001110100100001110",
7373 => "11101001111000100000010000100000",
7374 => "11111000111000101111000100010000",
7375 => "11111101110100101111101011110010",
7376 => "11111111111110101111010111101011",
7377 => "10010010111110010001000010101001",
7378 => "00010000111101011111000100100011",
7379 => "11101011110100110001100111010111",
7380 => "00001001110100011110010100010101",
7381 => "11100111111001110000001100010101",
7382 => "11111010111011001111000100001100",
7383 => "00000000110100111111111011111011",
7384 => "00001000111110111111111111110101",
7385 => "11000001000000100001101010111101",
7386 => "00000110000010101111110000001111",
7387 => "11110010110111100000111100001001",
7388 => "11110101111000111110101100010111",
7389 => "11110111111001110000100100001011",
7390 => "11110101111011001111100100010000",
7391 => "00011001111111000001010000001001",
7392 => "00011000000100110001011100000000",
7393 => "11111110000000110010010011111010",
7394 => "00000101000010010000011111111010",
7395 => "00001010000000110000001000010110",
7396 => "11101101111111110001101000100101",
7397 => "00001100000110100000001000000110",
7398 => "00001001000011110000110000011111",
7399 => "11110001000010011111100011110010",
7400 => "11110010111011101111101111110111",
7401 => "11110001111101011110110011110111",
7402 => "11111110111100101111100111111000",
7403 => "00000000000010111111101011111000",
7404 => "11111100111110001110100111111101",
7405 => "00000000111101100000010100000010",
7406 => "11110100111110001111111011110000",
7407 => "11111100111111001111010011110101",
7408 => "00001011111110111111100011110010",
7409 => "11110010111101111111101011110100",
7410 => "00000111111101011111011000000000",
7411 => "11111100111010111111101111111010",
7412 => "00000010111101111111010011111110",
7413 => "11110100111101011111010100000010",
7414 => "11111001111100101111101100000111",
7415 => "00000000111000001111110111111001",
7416 => "00001000111110110000010011111001",
7417 => "00000001111111100000100000000011",
7418 => "00000111000000110000001100010100",
7419 => "11110110110110010001000111101000",
7420 => "00001010000010011111011100001100",
7421 => "11101111111110011111111100000100",
7422 => "11111101111110111111111000000111",
7423 => "11111111111011011111100111110001",
7424 => "00001100111101110000111111111011",
7425 => "11111101111110110001000011111000",
7426 => "00010001111111100000000000011011",
7427 => "00000001111010000000100111100010",
7428 => "00010010000000010000000100010001",
7429 => "11110000111111001111010100010010",
7430 => "00000000111110001111101100010001",
7431 => "00001100111100110000110111111101",
7432 => "00000111000010000000000000000001",
7433 => "00001010000011000000101100000010",
7434 => "11111001000010010000101100001100",
7435 => "00001100111100111111000011011100",
7436 => "00001110000011100000101100001100",
7437 => "00001100000000111111010000000100",
7438 => "00000011000000100000001000001101",
7439 => "11111111111111100000001011110111",
7440 => "00001011111101011111110100000010",
7441 => "11111100000001010000100111110010",
7442 => "00000111000010010000011100000110",
7443 => "00000001000001000000000111101001",
7444 => "00001100000001111111101000001000",
7445 => "11111000000000011111010100000011",
7446 => "00000110111101111111110100001100",
7447 => "11110111111111101111101111111011",
7448 => "00001001111101010000101011110110",
7449 => "00010000111110110000101011111000",
7450 => "11111100000000010000000000000101",
7451 => "11111110000001110000111111101111",
7452 => "00010011000001001110110000000010",
7453 => "11111001111111001111010100001011",
7454 => "00000010111101101111101000001000",
7455 => "00000001111111101111100111110001",
7456 => "00001010111110100000110011101110",
7457 => "11100010111111010000101111011010",
7458 => "00010111111110011111101100000110",
7459 => "11110101111100110001000111011011",
7460 => "00010100111011101111011000001101",
7461 => "11111010111111111111111000011000",
7462 => "11111111111110001111001000001010",
7463 => "00000000111111001111110011111001",
7464 => "11111000111111111110001111110011",
7465 => "11110001000000010000001011101000",
7466 => "00101000111111011111110000001101",
7467 => "11111001110110010001010011000110",
7468 => "00010110111111001111110000001001",
7469 => "00000001111110011111110000011111",
7470 => "11111111000001001111110000000000",
7471 => "11111010111110011111010111110101",
7472 => "11110000000001011101110011110110",
7473 => "11001111111111111111100011001100",
7474 => "00001100000000111111011100010101",
7475 => "11110001111001010000010010101100",
7476 => "00001100111011011111111011111001",
7477 => "11110100111110111111110000010101",
7478 => "11111111111101011111010000000110",
7479 => "11111010111100001111010100000001",
7480 => "11111110111111111110010111110011",
7481 => "11100011111111010000010111100110",
7482 => "00010010111111001111000100011010",
7483 => "11110001110111000001100011010010",
7484 => "00001100111100111111011100001000",
7485 => "11111110111101000000011000001010",
7486 => "11111001111110101111101100001000",
7487 => "11111001111100011111010111110010",
7488 => "11100000000011001101011111101110",
7489 => "11100111000010101110000111110001",
7490 => "00001010000010011111101100000110",
7491 => "00000000110111010001010011101111",
7492 => "00000100111010001111011111111001",
7493 => "00000010111101110000100100000111",
7494 => "00000000111111101111111111101000",
7495 => "11111110111110101111101011111101",
7496 => "11111001111110001111110011110111",
7497 => "00000010111110010000101100000000",
7498 => "00001001111011001111100000000110",
7499 => "11101101111110010000110111101100",
7500 => "00000100111110110000010000010011",
7501 => "11100100000001000001000000000011",
7502 => "11110111111111101110111100000110",
7503 => "11110001000010001111100111100010",
7504 => "11111111111011111111111111101110",
7505 => "11100111111011011111010011110001",
7506 => "00000101111011111111010011111001",
7507 => "11110000000100101111001011111000",
7508 => "11100101111010111110101011111011",
7509 => "11111001111011001110000000000100",
7510 => "11110101111011101110111111110101",
7511 => "11110011111101011111010111101101",
7512 => "00010000111111010000001111110001",
7513 => "11110011111101010000111111110000",
7514 => "00001111111100001111001100000001",
7515 => "11110010110111100001100000001011",
7516 => "00010011111100101110110011110101",
7517 => "11100110111110010000010000001000",
7518 => "11111000111100001111010000001111",
7519 => "11111100111001111111110111110100",
7520 => "00011001111101110001100011110111",
7521 => "11101101111110110001011011110000",
7522 => "00011001111110111111100000001101",
7523 => "11111010111001000011001000000101",
7524 => "00100000111101001111100100001001",
7525 => "11101101000000000001010000001001",
7526 => "11111101111100101111111000010111",
7527 => "11111111111011000000000011110010",
7528 => "00001101111110010001000011110000",
7529 => "11101101111110110001110111101010",
7530 => "00110001000000101111011000011011",
7531 => "11101001110111110010111111101010",
7532 => "00011100111110111110111000010010",
7533 => "11101011111100000000000000010001",
7534 => "11111010111100011111101000010101",
7535 => "00001001111000100000110011101000",
7536 => "00000100000001100000010011111000",
7537 => "11101001111101110001010111101111",
7538 => "00100111000000001111101000011001",
7539 => "00000000111001010000110011100000",
7540 => "00011001111101000000110100001101",
7541 => "11111001000001111111001100011110",
7542 => "11111011111111111111100000001110",
7543 => "00000110111011110000011011101011",
7544 => "00000001000000000000010111111100",
7545 => "11110000111111100000011011100101",
7546 => "00100000111111101111111000001010",
7547 => "11111011111110000001001111110101",
7548 => "00001111111110100000010000000111",
7549 => "11110111111111011110110100001100",
7550 => "11111001111110100000000100000001",
7551 => "11110100000100001110111111110011",
7552 => "11111101111011010000100111110100",
7553 => "00000011111101110000011111111000",
7554 => "00000000111101101111100000000000",
7555 => "11110101000010110000111011111001",
7556 => "00001011000000001110101100000011",
7557 => "11111001111100111111110000010001",
7558 => "11110001111011111111011100000011",
7559 => "11110101000000101111100011110011",
7560 => "11110001111100001111101111111010",
7561 => "11111100111100101111101111111010",
7562 => "00010111111100011111100100000000",
7563 => "11110011111100110000100011101011",
7564 => "00001000111111101111011011111111",
7565 => "11110010111100101111110000011010",
7566 => "11110110111101111111001111111000",
7567 => "11111110000000100000000111110010",
7568 => "11101111111111101101110111111111",
7569 => "11110110111110001111010011111100",
7570 => "00011111111101101111101000001111",
7571 => "11111100111011000000000011001101",
7572 => "00001011111110111111111100000001",
7573 => "00000001111110111111111100010101",
7574 => "11111100000001010000001011111001",
7575 => "11111010000000111111110111111111",
7576 => "11100111111111101101010100000010",
7577 => "11110101111110111111000011110111",
7578 => "00011011111110000000000000001111",
7579 => "11110101111101101111110111010011",
7580 => "00000101111100111111011011111000",
7581 => "11110000000001101111101000010100",
7582 => "00000000000000111111111011111110",
7583 => "11111111000000011111100100001100",
7584 => "11110001111110111101110000000010",
7585 => "00000011000000111111101100010000",
7586 => "11111100111110101111111100010011",
7587 => "11111000111101001111111111100010",
7588 => "00000000111110011111100100000100",
7589 => "00000010000000000000010000000111",
7590 => "11111110000000110000001111111100",
7591 => "11111010000000011111101100001010",
7592 => "11110100000000011110111000000111",
7593 => "00000100111101101111000100011000",
7594 => "11111101111110101111011000010000",
7595 => "00000101111101100000000111100000",
7596 => "11110111000001110000001111110110",
7597 => "00001010111111000000011111111101",
7598 => "11110100000000010000101111110100",
7599 => "11111011000000111111001111110100",
7600 => "00001000111101100000110011111010",
7601 => "00000000111100100000000100000011",
7602 => "00000000000001011111101111111100",
7603 => "11100101000000011111000100001001",
7604 => "11111001000000001110000011110010",
7605 => "11101100111011011111100000000000",
7606 => "11110110111111011111011111110101",
7607 => "11101110111111111111100111101111",
7608 => "11111010111000011111010111100101",
7609 => "11100010111011011110111111110000",
7610 => "11111111111100111110110111111000",
7611 => "11111010000001100000110000001011",
7612 => "00001000111000001111001111101100",
7613 => "11110100111101110000101100000011",
7614 => "11101110111011011111011011111010",
7615 => "11111011111110101111000011111110",
7616 => "00010110000001000000010111111101",
7617 => "11111110000010010000010111111001",
7618 => "00001100111111011111100000000000",
7619 => "11111000111011110000011100010000",
7620 => "00001011111110111111010011111011",
7621 => "11110000111101100000110000000101",
7622 => "11111110111110001111011000001111",
7623 => "11111111111100111111100100000000",
7624 => "00000110000000100001001011111100",
7625 => "11110010000011010000000011110011",
7626 => "11111110000000101111100111110111",
7627 => "00000000111001000001011000001111",
7628 => "00000110111111111111111111111000",
7629 => "00001110111111110000111000001000",
7630 => "11111111000000000000000100000011",
7631 => "11101100111011011110111011111000",
7632 => "00001011111100010000100011110110",
7633 => "11101111111101000001010011101000",
7634 => "00100110111110101111110100011001",
7635 => "11101100110111100001110000000110",
7636 => "00010111111101101110010100000110",
7637 => "11101011111011100000000100011000",
7638 => "11111001111010111111011000010010",
7639 => "11110011110100001111101011101111",
7640 => "00000001111111100001000111101100",
7641 => "11100111111100000001100011101010",
7642 => "00101111111101111111100100100010",
7643 => "11110100110100100010010000000011",
7644 => "00001111111100101111100000001111",
7645 => "11101100111100100000100100011001",
7646 => "11111100111010001111000000010010",
7647 => "11101110111011101111111011110001",
7648 => "11111001111110010000010111110010",
7649 => "11100101111110010000011111010100",
7650 => "00100001111101001111011000001001",
7651 => "11111001111100000001001100001011",
7652 => "00001010111100101111010011111110",
7653 => "11111010111101010000010100011001",
7654 => "11110111111011111111110100000001",
7655 => "11111000111110111111101011111000",
7656 => "11110001111110111111111011111000",
7657 => "00000110111101011111001011111101",
7658 => "00001001111100111111101100000101",
7659 => "11111110111110110000110100000001",
7660 => "11111111000000111111110011110000",
7661 => "11111001111111100000010000001000",
7662 => "11110110111111111111111111111101",
7663 => "11111001000000111111100011111111",
7664 => "00000001111111111111111011111101",
7665 => "11111110111111101111100111111110",
7666 => "00000001111110110000000000000000",
7667 => "11111010111101101111111111101111",
7668 => "11111110111111111111101111111110",
7669 => "11111110111111101111111100011010",
7670 => "00000000111110100000000100000000",
7671 => "11111101000001011111110000000000",
7672 => "11111000111101101110011000000101",
7673 => "11111111111111101110111000000010",
7674 => "00011000111111100000000000000010",
7675 => "11110100111101011111111111101000",
7676 => "11111111000000101111101111111001",
7677 => "11111000000000000000100000010000",
7678 => "11111110000001011111111111111111",
7679 => "00000000111111001111111100000100",
7680 => "11101001000001111110101000000011",
7681 => "11111111000000011110000100000100",
7682 => "00010001000001010000011000000010",
7683 => "00000010111110011111110011101010",
7684 => "11111000111111000000010011111011",
7685 => "11111110111111001111100000001101",
7686 => "00000000111111110000011011101010",
7687 => "00000011000000001111111100001110",
7688 => "11111000111111111111000100000000",
7689 => "11111101000010011111011000001110",
7690 => "11111110000001110000010000000011",
7691 => "11111110111111001110101111110100",
7692 => "11110011111111001111110111111100",
7693 => "11111100000000011111011100001001",
7694 => "11111111000001010000010111110110",
7695 => "11111100000000110000011011111001",
7696 => "11101100111110111111010111111111",
7697 => "11110111000000111110010011101100",
7698 => "00000000111110000000010011101010",
7699 => "00000011111111101110110111101101",
7700 => "11111011000000000000101011011110",
7701 => "00000110000010101111001000000100",
7702 => "00000100111111110000000011100101",
7703 => "11111001111111101111101011111101",
7704 => "11110110111101001111101000000000",
7705 => "00000111111110001110111100000110",
7706 => "00000011111101011111110111110011",
7707 => "11111000111101000000101100000011",
7708 => "00000011000000011111100111110111",
7709 => "11110000000001000000100100000101",
7710 => "11111001111110111111101011110111",
7711 => "11111000111111011111011011111101",
7712 => "00000010000001010000010111111111",
7713 => "11101100000001101111110011101101",
7714 => "00000010111101011111100111111000",
7715 => "00000000000000100000100011111111",
7716 => "00000110111010010000000111110111",
7717 => "00000001000000000000000011111110",
7718 => "00000001111110111111111111110110",
7719 => "00001010000100001111110111111100",
7720 => "00000100000000100000100111111101",
7721 => "11111101111101100000011011110111",
7722 => "00010000000000011111110000000001",
7723 => "11111000111101010000011100000000",
7724 => "00000011111101100000010100000001",
7725 => "11111000111111111111110000001011",
7726 => "11111010111110111111111000000000",
7727 => "00000101111101010000000111111111",
7728 => "00001010000000100001100111111011",
7729 => "11111000111111100001000011110001",
7730 => "00010100111110111111011100001101",
7731 => "00001000111101000001111100001100",
7732 => "00010100111101100000011100000101",
7733 => "00001010000000100000011000001010",
7734 => "11111101111111110000000100001110",
7735 => "11111110111011001111010100000110",
7736 => "00000110111111010001000111111010",
7737 => "11110110111111110000110111101111",
7738 => "00010101111110001111111100000111",
7739 => "11110101111001100001110000001010",
7740 => "00010001111111011111100100000000",
7741 => "11101110000000000000110100001001",
7742 => "00000011000000101111011000001011",
7743 => "11110010110111001111000000000100",
7744 => "00000010111101110000110011111010",
7745 => "11110100111111100000000111101110",
7746 => "00010110111110111111101000000010",
7747 => "11110101110101000001001000001010",
7748 => "00000100111110001110110011111111",
7749 => "11110101111101000000010000011000",
7750 => "00000000111101011111111000000100",
7751 => "11101010111001111111100000000100",
7752 => "11111001000000010000110011111011",
7753 => "11111010111110111111101111101110",
7754 => "00010000111111001111111011110110",
7755 => "11111101110110110001001000001011",
7756 => "00001101111111001111000111110111",
7757 => "00000001111111100000100100011001",
7758 => "11111011111110001111101000000010",
7759 => "11110001111110011111011000001011",
7760 => "00000000111100100000100111111111",
7761 => "11111111000000000000010011111100",
7762 => "00001110111110101111100100000010",
7763 => "11111000111011110000101000000011",
7764 => "00001011111111111111000011110101",
7765 => "00000001111110010000110100010000",
7766 => "11111100111110101111101000000111",
7767 => "11111101111100011111011100000110",
7768 => "11110111111101000000000100010000",
7769 => "00000000111111101111101000000011",
7770 => "00001000111111110000000011111001",
7771 => "11111111111110000000001100001011",
7772 => "11101101000000011111110111110001",
7773 => "11110111000000110001000000010100",
7774 => "11111010000001100000010011111000",
7775 => "11111101111111110000001100000100",
7776 => "00000010111110110000001000000011",
7777 => "00000101111111001111011100000110",
7778 => "00001011111111110000101111111110",
7779 => "00000010111111110000000100001000",
7780 => "11110110111111110000000011110100",
7781 => "11111110000011100000000100000011",
7782 => "11111111000001100000100111110011",
7783 => "00000111000001000000001000000000",
7784 => "11111001000000001111111100000111",
7785 => "00001011111110111111101000000110",
7786 => "00010011000000100000010111111100",
7787 => "00000000000000011111001100000110",
7788 => "11101101000001010000001111111110",
7789 => "00000101000011100000011100001111",
7790 => "11111111000010000000101011110011",
7791 => "00000011111111100000001000000001",
7792 => "11110001111111011110111011111110",
7793 => "00001001111101011110010000001011",
7794 => "11111110111100010000001100000100",
7795 => "00000101000000001111000011111011",
7796 => "11101001000010010000001011110000",
7797 => "00000100000000101111100100000101",
7798 => "00000110000010110000011111101010",
7799 => "00000000000010000000110000000111",
7800 => "11101100000010011110110011111110",
7801 => "00001011111101111110001100001110",
7802 => "00000001111111100000001011111101",
7803 => "00001111000000011110111011100011",
7804 => "11111111000001000000110011101011",
7805 => "00001010111110111110110111111101",
7806 => "00001001000011010000001011101101",
7807 => "11111111000001000000000011111111",
7808 => "11100100111100111110011000000000",
7809 => "00000111111110111110011100000111",
7810 => "00000001111001111111111011111110",
7811 => "00001011111110110000101011110011",
7812 => "00000110000000001111000011110110",
7813 => "00010000111101110000001100000000",
7814 => "00000100111111100000011111111001",
7815 => "11110111000000010000000111111011",
7816 => "11110011111011000000011111111110",
7817 => "11110100111110101111010111111011",
7818 => "00000100111101011111101111111110",
7819 => "11111110000001101111111000000101",
7820 => "11111001111101111110101011111010",
7821 => "00000000111101101111011000000000",
7822 => "11111010111110011111111011101111",
7823 => "11111001000011010000000100000001",
7824 => "11111000111111011111001111111010",
7825 => "00000001111110101111011000000100",
7826 => "00000110111100101111110111111011",
7827 => "00001000111101110000100100001000",
7828 => "00000110000001100000011011111110",
7829 => "11111101000000100000101100000110",
7830 => "11111001000000000000001111110111",
7831 => "00000001111011010000001000000000",
7832 => "11111110111111110000001111111101",
7833 => "11111101111110011111100111110101",
7834 => "00000100000000111111110111110110",
7835 => "11111100000010110010011100011100",
7836 => "00001011111110110000000111111011",
7837 => "00000110000000000001001100000011",
7838 => "11111110111110110000000011111010",
7839 => "00000010111001100000000100000101",
7840 => "00000110000001110000001100000010",
7841 => "00000101000001100000110000001010",
7842 => "00010110000000000000000000000110",
7843 => "11110110000010100001010000101010",
7844 => "00000010000001111111110100000111",
7845 => "11110000000000110001001000000101",
7846 => "00000000000000110000001100001000",
7847 => "00000101110111000000011000001101",
7848 => "00000011000001110000001000000100",
7849 => "00000000000011010000010111111101",
7850 => "00000111000001100000010011111101",
7851 => "00000001111100010001011000011001",
7852 => "00000111000000100000011000000001",
7853 => "11111101000001000000111000001101",
7854 => "00001000000001000000101100000101",
7855 => "00000000110100110000000000001010",
7856 => "00001010000001000000011000000110",
7857 => "11111100000100100000000011110101",
7858 => "11110011000010100000101011110100",
7859 => "00000101111011000001001111111001",
7860 => "00000011111111101111110100000010",
7861 => "00000000111111110000100100001000",
7862 => "00001010000000100000101000000001",
7863 => "11111110111000100001000000010000",
7864 => "00000111111111100000111000001001",
7865 => "11111110000001110000010011111010",
7866 => "11101111000011100000011011110000",
7867 => "00001010111101010000011100000001",
7868 => "11110111000000001111100011111110",
7869 => "00001010000001100000100000010010",
7870 => "00000010111111100000100100001100",
7871 => "00001010111101000000010000000111",
7872 => "11111110000000110000011000001100",
7873 => "11111101000010011111101111111100",
7874 => "11110110000010110000110011110000",
7875 => "00000001000001000000011100000110",
7876 => "11110011000000000000000011111000",
7877 => "00000001000010000000100000000101",
7878 => "00000110000000100000010111111100",
7879 => "00000011111101100000000000001110",
7880 => "11111101111110000000101000001011",
7881 => "11111011000000111111101111111111",
7882 => "11110000000001110000101111010111",
7883 => "00000001000000101111110100010100",
7884 => "11100010000000100000001011110001",
7885 => "00000101000010110000001100000111",
7886 => "00001100000000100000000011110111",
7887 => "11111101111111001111011100000111",
7888 => "11111011111100100000011100000110",
7889 => "00000000000000011111100000000111",
7890 => "11111011111110000000001111010011",
7891 => "00000101000001011111110100011000",
7892 => "11100111111111111110101111101111",
7893 => "00001100000000110000001000000010",
7894 => "00000100000000010000110111110010",
7895 => "00000011000000010000010000001111",
7896 => "00000101111110010000000100001010",
7897 => "00011000000001111111100100010101",
7898 => "11110111000000100000010111110001",
7899 => "11111100000001011110111100010111",
7900 => "11100010000011011111011011111011",
7901 => "00000010000001110000101000000010",
7902 => "11111111000010000000101011111100",
7903 => "00000011000010100000011000000000",
7904 => "00000000000001010000101000001011",
7905 => "00001010000010001111011100010001",
7906 => "11111100000001000000111011110111",
7907 => "00001001000001101101111000001110",
7908 => "11110011000100000000010011111101",
7909 => "00000110000011001101100100000011",
7910 => "00001011000101010000100011111101",
7911 => "00000110000100100000101011111000",
7912 => "11111100000010101111100100000001",
7913 => "00000100000001011111010100000100",
7914 => "00000001000011100000010011111010",
7915 => "00010010000010110000000111110100",
7916 => "00011001111101110000010111111011",
7917 => "00010101000001101111101011111111",
7918 => "00001000000000010000111011111011",
7919 => "11111101000000101111111100000100",
7920 => "00000011000001010000000000000011",
7921 => "00001001111111101111010100001110",
7922 => "00000000111111110000000100000010",
7923 => "11111100000010010000001100000011",
7924 => "11111010000001110000010000000010",
7925 => "00000000000001100000011000000101",
7926 => "00000010000010001111111100000001",
7927 => "00000000000010111111110111111010",
7928 => "00000010000010100000000100001000",
7929 => "11111010000001110000000011111001",
7930 => "00000011000010001111111000000111",
7931 => "11111011111111101111101011111100",
7932 => "00001001111111100000000100000000",
7933 => "00001000111101100000100000000100",
7934 => "00000011111110010000000100000110",
7935 => "11111111000001011111110111111011",
7936 => "11111101000000101111101011111110",
7937 => "11111011000010111111011111111010",
7938 => "00000011000010111111101100000010",
7939 => "11111010111111000001001100000100",
7940 => "00011001111111011111111000000010",
7941 => "11111001000000100000000000000001",
7942 => "00000101111100101111111111111111",
7943 => "00000101111001011111100100001001",
7944 => "00001001000010001111110000000001",
7945 => "00000110000010000000010100001010",
7946 => "11111110000001010000010000001011",
7947 => "11111101111010000001110100010100",
7948 => "00010011000001100000010000000111",
7949 => "11111100000010100001011011111101",
7950 => "00000001000001101111110000001100",
7951 => "00000010111011101111110100000000",
7952 => "00000110000010111111110100010000",
7953 => "11101110000001000000010011110100",
7954 => "00001000000010100000001111111111",
7955 => "00000101111110000010011011111010",
7956 => "00010111111101000000011100001001",
7957 => "00000010000000100001011100000111",
7958 => "00000111111111101111110100000100",
7959 => "00001011111001100000101100001110",
7960 => "00001100000011000000011100000000",
7961 => "11110110000000000000100111101111",
7962 => "00001000000010000000100111111111",
7963 => "11111011111110110010001000101001",
7964 => "00001010111111100000110000000111",
7965 => "11111001000001000001010000000110",
7966 => "00000100000010000000011100000110",
7967 => "00010001111011000000110000010010",
7968 => "00001100111110110000101100000101",
7969 => "11111001000010100000101011110111",
7970 => "11110111000010010000001111110010",
7971 => "00001011000001110001110000100111",
7972 => "11110101111110010000011100000100",
7973 => "11111111000011100001101000001101",
7974 => "00000100000100100000101000000111",
7975 => "00000101111100010000010100001100",
7976 => "00000101111110000000000100001101",
7977 => "00001111000001000000000100000010",
7978 => "11101011111110110000010011101101",
7979 => "11111111000011000000001000101001",
7980 => "11010100000001011111100011111110",
7981 => "00000101000011000000110111111101",
7982 => "00000010000010010000100011111101",
7983 => "11111100111101011111101000001100",
7984 => "00000101111110100000010000000111",
7985 => "11110000111111001111111011111010",
7986 => "11110110000000100000001011011100",
7987 => "11111111000010100000001000001001",
7988 => "11001010111100101111011011110110",
7989 => "11111100000000100001000100000111",
7990 => "00000110000000110000101011110110",
7991 => "11111111111111000000001100001001",
7992 => "11111101111110000000100100001100",
7993 => "11111110111100001111110000001011",
7994 => "11111011111110110000010011100100",
7995 => "00000101000001101111000000001111",
7996 => "11011010000000001111011111110101",
7997 => "00001000111111101111011111111100",
7998 => "00000010000001100000010011110101",
7999 => "11111111111111000000010100001001",
8000 => "00000001000000000000001000000011",
8001 => "00001001111110111111110100001111",
8002 => "00000010000000100000000011110011",
8003 => "11110011000001011110110000010110",
8004 => "11100010000010111110111111111111",
8005 => "11111001111100110000111000000001",
8006 => "11111101000000110000100011111011",
8007 => "00001101111111100001100000000000",
8008 => "00000101000001111111111100001100",
8009 => "00010000000001010000001100010110",
8010 => "11111100000000010000010100001001",
8011 => "00000100000001001111001011111111",
8012 => "11111001000001001111111100010001",
8013 => "11111101000010011110111011111100",
8014 => "00000110000011010000100100000011",
8015 => "00001001000101100000101100000011",
8016 => "00001001000011100000111100000000",
8017 => "00001101111111110000100011111111",
8018 => "00000010000010000000001000000111",
8019 => "00001000000101101111101000000100",
8020 => "00001110111111010000101000010000",
8021 => "00000111000100000000110100000000",
8022 => "00000110000011110000001100001111",
8023 => "11111011000001000000001000000011",
8024 => "00000100111111111111100100000101",
8025 => "00001011000000011111101100001000",
8026 => "00000001000000110000001011111111",
8027 => "00000001000001110000000100000100",
8028 => "11111010000010000000000100001100",
8029 => "00000010000000110000011000000110",
8030 => "00000100000010011111111100001101",
8031 => "00000100000100000000010111111011",
8032 => "11110101000010001111010111111000",
8033 => "11100011000000111111001011110011",
8034 => "00000010000000101111101111111100",
8035 => "11111110000010001111110011111110",
8036 => "11111001111010001111101111101001",
8037 => "00000011000000011111000000000101",
8038 => "11111111111110001111100111101000",
8039 => "00000100111011010000000111101010",
8040 => "11111010111011011111110011111110",
8041 => "11100110111011001111110111110100",
8042 => "00000001111011111111011100000010",
8043 => "11111000111010001111111011110010",
8044 => "00000011111110011110111011111011",
8045 => "11110111111011111111100000000001",
8046 => "11110011111101011111110111111001",
8047 => "00001001111000010000101011110011",
8048 => "11111101111110010000010111111001",
8049 => "11110000111100010000101111111000",
8050 => "00000100000000110000000000000100",
8051 => "11111011111100011111100111101110",
8052 => "11110100111011011111110100000101",
8053 => "11111101111111011111000100000001",
8054 => "11111010000001000000000111111110",
8055 => "00001101111010100000110000000000",
8056 => "00000010000000010000001011111101",
8057 => "11111000111101000000011111111001",
8058 => "11111011000000100000010000001001",
8059 => "00000011000000111111110100001000",
8060 => "11101011111110100001100100000111",
8061 => "11111100000100101110101100000011",
8062 => "11111010000010101111110111111011",
8063 => "11111101111010001111010100001011",
8064 => "00001011000010100000100000001111",
8065 => "11110010111110110000101100000010",
8066 => "00000011111110000000010100001100",
8067 => "00000101111011100001000011111011",
8068 => "00001100111111111111101100001100",
8069 => "11110110111101000001011011111011",
8070 => "00000001111101110000010100001110",
8071 => "00001000111101010000001100000000",
8072 => "00001101000000100000100100000100",
8073 => "11101011000001010000111111110000",
8074 => "11111000000010010000011000000101",
8075 => "11110110000001100001000100001000",
8076 => "11111100111110010000001100001000",
8077 => "11111110000001100000101000000000",
8078 => "00000100111110010000000000010000",
8079 => "00001000111100110000001100001011",
8080 => "00010010000010000000111000010010",
8081 => "11111101000101010000110011111110",
8082 => "11110110000011110000011000000011",
8083 => "11111010000001110000111100010000",
8084 => "11011111000000111111100100010000",
8085 => "11111011111111110010001011111111",
8086 => "00000110000000110000010100010010",
8087 => "00010000000000000000011111111001",
8088 => "00010100000001100000110100000111",
8089 => "11101100000100110000110011101011",
8090 => "11110110000100110000011000000001",
8091 => "11111111000011000000011100000101",
8092 => "11001010111100110000010100001000",
8093 => "00000010000010110001000000000010",
8094 => "00000111000000111111111100001101",
8095 => "11111100000011001111110011111110",
8096 => "00010000000001000000101100000001",
8097 => "11110100000101010000001111111000",
8098 => "00000001000100010000000111111001",
8099 => "00000001000100011111110100010111",
8100 => "11101101111101111111011111111111",
8101 => "00000011000001000001010000000110",
8102 => "11111011111111001111111000000101",
8103 => "11111001111101011111110000000101",
8104 => "00001110111111000000011000001010",
8105 => "00001100000001101111111000001101",
8106 => "00000000000010010000001011111101",
8107 => "11110111111110011111010100001110",
8108 => "11101011000010111110101100000111",
8109 => "11110101000000010000100000000110",
8110 => "00000011000001110000011000000011",
8111 => "00000010000010100000010100000100",
8112 => "00001001000011110000101100000010",
8113 => "00010011000011010000011000010001",
8114 => "00000100000011100000010000001000",
8115 => "11111101000001101111010011111111",
8116 => "11111001000000100000000100001100",
8117 => "00000000000001101110101000000001",
8118 => "00000111000000110000010000001100",
8119 => "00000100000101000000000000000011",
8120 => "00010011000001000001000011111110",
8121 => "00001011111111000001000000000111",
8122 => "11111111000010100000010111111111",
8123 => "00000000000101011111110000010000",
8124 => "00001110111111101111110000001000",
8125 => "11111111111111111111101100000100",
8126 => "00000111111111100000010000000100",
8127 => "00000000000000000000000000000000",
8128 => "00000000000000000000000000000000",
8129 => "00000000000000000000000000000000",
8130 => "00000001111111101111110100000000",
8131 => "00000000000000011111110111111110",
8132 => "11110100111111010000010011111110",
8133 => "00000000111111100000001111111101",
8134 => "11111100111110100000010011111110",
8135 => "11111001111111000000001100000001",
8136 => "11111101000000000000001000000010",
8137 => "00000000111111010000001000000001",
8138 => "11111101111101110000001100000011",
8139 => "00000000000001010000001000000001",
8140 => "00000111000000110000010011111110",
8141 => "00000100000000100000001111111111",
8142 => "00000101111110010000000000000000",
8143 => "11111100000001110000011000000011",
8144 => "11111110000000000000000000000100",
8145 => "00000110000000011111111100000011",
8146 => "00001001111111100000011100010101",
8147 => "00000001000000101111111100001101",
8148 => "00010011000011100000100100001110",
8149 => "11111111000010100000111000000011",
8150 => "00011011111110110001000000001011",
8151 => "00010010000001110001010000000100",
8152 => "00000111000101010001101000000011",
8153 => "00001000000010100000111100001010",
8154 => "00010001000100100000101100001111",
8155 => "11111000000011001111110100000110",
8156 => "00010010000010010000111100001110",
8157 => "00000001000100000000101100000010",
8158 => "00001100000101100001111000010001",
8159 => "00011100000001000001010100001101",
8160 => "00001101000001110000111111111100",
8161 => "00000111000001000000100100000111",
8162 => "00010100000110011111100000000110",
8163 => "11111101000010011111111000001010",
8164 => "00001111111111010000010000001110",
8165 => "00000100000100000000100011111101",
8166 => "00000111001000110000000100000111",
8167 => "00000101000001101111111000001100",
8168 => "00010011000000010000100000000010",
8169 => "00001011000001010001010000000100",
8170 => "00000011000100011111011100000000",
8171 => "11110111111111011111110000001011",
8172 => "00011010000001111111011100010111",
8173 => "00000011000001100000110100000001",
8174 => "00010001000101010000001100001010",
8175 => "00001000000001100000101111110110",
8176 => "00001101000001000000011100000000",
8177 => "00001000000000110001000011111111",
8178 => "00001111000110101111111100001110",
8179 => "00001011001000000000001000001011",
8180 => "00010101000001001111011100010110",
8181 => "00000101000101010000010011111011",
8182 => "00010110000111110000110100001000",
8183 => "00001101000110100000111111111110",
8184 => "00000111000101100001011100000000",
8185 => "00000001000011100000000011111100",
8186 => "00000100000100101111011100000110",
8187 => "00010010000100000000001000001010",
8188 => "00000111000010111111111000000110",
8189 => "00000110000000110000010111111110",
8190 => "00000010000110110000010011110111",
8191 => "00000011000011010000001000000000",
8192 => "00001100111111110000010111111010",
8193 => "00001000000000110000101100000010",
8194 => "00001001000000001111110011111101",
8195 => "00011110000111100000101100000110",
8196 => "00010101000110010001100000000111",
8197 => "11111111000101100000100100000111",
8198 => "00000110000110011111110000000100",
8199 => "11111111000011100001010000010001",
8200 => "11111111111111011111110111111100",
8201 => "00001010000000100000001100011001",
8202 => "00000010000010100000001000001110",
8203 => "00010010000111000000100100000111",
8204 => "00011111000101110001100000010101",
8205 => "00000100000011010000011100000011",
8206 => "11111111000111000000111100001010",
8207 => "00001111000101100001010100010101",
8208 => "00000111000011100000011011111100",
8209 => "00001111000001000000110100000100",
8210 => "00001011000010000000010100001011",
8211 => "00010000000101000000010100000110",
8212 => "00010100000110110000110000000111",
8213 => "11111111000011010000101000000010",
8214 => "00001110000111000001000100001011",
8215 => "00010010000011100000010000001010",
8216 => "00000110000010000000100000000001",
8217 => "00001101000001110000011000000111",
8218 => "00001011000101010000110100001010",
8219 => "00001011000000010000100000001010",
8220 => "00011010000010100000000000001101",
8221 => "00001000000010110000110000000010",
8222 => "00001100000100000001001100001010",
8223 => "00010110000001100001000000000001",
8224 => "00010110000010100001100111111101",
8225 => "00001101000010100001000000000011",
8226 => "00000101000011010000011000000101",
8227 => "00000000000000000000000100000001",
8228 => "00000111111111010000010000000110",
8229 => "11111111000000000000001100000000",
8230 => "11111101000011010000111000000110",
8231 => "00001111000001010000001011111101",
8232 => "00000111000000100000111100000011",
8233 => "00000101000000110000010000000001",
8234 => "00000011111110110000010011111010",
8235 => "11101111111111100000000000000010",
8236 => "11100110111110101111101011110011",
8237 => "00000011111111101111110000000000",
8238 => "11110100111101101111111011111110",
8239 => "11111010111100011111110011110111",
8240 => "11110101111110111111110000000001",
8241 => "00000010111111101111111111111000",
8242 => "11111110111010101111111000001001",
8243 => "11101110000001101111100111111110",
8244 => "00001101111111101111100000010001",
8245 => "11111111000001001111110100000010",
8246 => "00000101111011000000111000001110",
8247 => "00000101000011000000100100001111",
8248 => "00000100000011100001000111111110",
8249 => "11111111000011000000011011111110",
8250 => "00000011000101010000101000000101",
8251 => "11111100000000110000001000000011",
8252 => "00001110000010000000101000001101",
8253 => "00000001000001010000011000010010",
8254 => "00010010000011010001001100000001",
8255 => "00010001000001000000011100010110",
8256 => "00010111111101110000101111111110",
8257 => "00000100111111110000010011111110",
8258 => "00000000000011000000010000000011",
8259 => "11100100000010111111010100001010",
8260 => "00001101000000011110011000001001",
8261 => "11111100000000111111111111111110",
8262 => "00010100001000010000100000000011",
8263 => "00000011000010100001000100000111",
8264 => "00001100000010110000111111111011",
8265 => "00000001000010100000111111101100",
8266 => "11110111001000111111100100001000",
8267 => "11101011000000011111100000000011",
8268 => "00000111000001111101110000000111",
8269 => "11111110111101110000001011101011",
8270 => "00001101001001011111100111111101",
8271 => "00000100000010001111111011101101",
8272 => "00010111000000010000011011111001",
8273 => "11111110000001110000011011100110",
8274 => "11111110001000111111101011111101",
8275 => "11101000111101001111110100000001",
8276 => "00000111111110001101100000000111",
8277 => "00001001111101101111110011100001",
8278 => "11111001001010101110100011110111",
8279 => "11110100000010001111001011011101",
8280 => "00001001111110011111101000000010",
8281 => "11111001111111110000101111100011",
8282 => "11111100000011010000101111110111",
8283 => "11110100111011101111111100000100",
8284 => "00001001111110011101101100001100",
8285 => "00000000111100110000001111101111",
8286 => "00000011000100111111000100000100",
8287 => "11110111111111100000011011100101",
8288 => "00000111000000101111010100000110",
8289 => "11111010000000101111111111011100",
8290 => "11111011000001110000100011111110",
8291 => "11111100111010100000101011111101",
8292 => "00000000111110101111100100001000",
8293 => "00000101111011101111110011101001",
8294 => "00000001000100001111010000000100",
8295 => "11111001111111111111011111100011",
8296 => "00000001000000010000000100000011",
8297 => "11110100000001000000011111110110",
8298 => "11111110111111100000001011111110",
8299 => "11110111111100010000000100001001",
8300 => "00000011111100101110111000001000",
8301 => "11111001111110010000011011111110",
8302 => "00000001000000011111000000001100",
8303 => "11110110000011011111011111110000",
8304 => "11111010111111111111101011110010",
8305 => "11110110000000110000000011101100",
8306 => "00001100111111110000101000000100",
8307 => "11110011111101111111010100001100",
8308 => "00010010000000001110111000010010",
8309 => "11111010000000100000111000000001",
8310 => "00000011111111101111011000001001",
8311 => "11110111000101101111110111110100",
8312 => "11111111000100100000000111110101",
8313 => "00000101000011000000011011110101",
8314 => "00001010000001111111110100000010",
8315 => "11111110000001100000011000000110",
8316 => "11111111000001110000110000000001",
8317 => "11111111000001010001000000000001",
8318 => "00000010000000110000001000000011",
8319 => "00001010000001100000011000000101",
8320 => "00000011000001111111111000000000",
8321 => "00000111000000101111111100000101",
8322 => "00001010000001000000011000000001",
8323 => "00001010000000010000000100000100",
8324 => "00010001000010101111110100001100",
8325 => "11111101000001010000100000000001",
8326 => "00000010000001010000001100000101",
8327 => "00001011000010010000000111110100",
8328 => "11111110000010011111111011111100",
8329 => "00000101000000110000100011111011",
8330 => "00000011000001000000010000000101",
8331 => "00000011000000000000010111111111",
8332 => "00000110000001111111000000000000",
8333 => "00000001000000011111111100000011",
8334 => "00000110000001110000101100001000",
8335 => "00000111000000000000000111110101",
8336 => "11111110000000010000101100000011",
8337 => "11111101000000000000000011111010",
8338 => "11110110000000001111111011111001",
8339 => "11110000111110001111101011111011",
8340 => "11100100111110001110110111110100",
8341 => "00000010111110111111100011111111",
8342 => "00000000111100100000001000000001",
8343 => "00000010111011111111011111111000",
8344 => "11111101111111000000000000000010",
8345 => "11111011111110111111101111101101",
8346 => "11111100111010111111111000000101",
8347 => "11111010000001011111101000000000",
8348 => "00001110000000101111101100001110",
8349 => "11111011000000000000000100001111",
8350 => "00001010111010110000010000000010",
8351 => "00000100000001010000101000001100",
8352 => "00001000000000000000101111111110",
8353 => "00000100000010001111111011111000",
8354 => "11111111000110110000000111111000",
8355 => "11100111111110110000000100000000",
8356 => "00010001111110111110110100001010",
8357 => "11111111111110010000011000001010",
8358 => "00000111000110011111100011110101",
8359 => "00001000000001111111111100001010",
8360 => "00010001111111111111001000000010",
8361 => "00000001111111101111111011110001",
8362 => "11111111000011100000000000000000",
8363 => "11100110111110011111001100000100",
8364 => "00001111000000001101110000010011",
8365 => "11110111000000000000010000000101",
8366 => "00001000000111001101011011111011",
8367 => "11101011000010100000001111111100",
8368 => "00001001111110101111101111111100",
8369 => "11111111000000100000011011100101",
8370 => "11110110000101110000010011110111",
8371 => "11101011111100010000010000000100",
8372 => "00000001111110001100101000000100",
8373 => "11110010111101000000001111011011",
8374 => "00000101000110111101101011110011",
8375 => "11101100111111011111101011010011",
8376 => "00001010111111011110100100000011",
8377 => "11111111111111111111110111011010",
8378 => "11110011001001111111011011110111",
8379 => "11101010111100011110111011111111",
8380 => "00000110000000011100011111111111",
8381 => "11110111111010011111011111010110",
8382 => "11111011000110111101111011111011",
8383 => "11011011000000101110111111011000",
8384 => "00001011111101101110110100001001",
8385 => "11111100111110101111110111011010",
8386 => "11110011000010001111011100000011",
8387 => "11111000111101001111110000000001",
8388 => "00001000111110101110010100001001",
8389 => "11100010111101110000000011011111",
8390 => "11110111000100101101101000000010",
8391 => "11001100000000101111010111100010",
8392 => "11111000111101011111010000001111",
8393 => "11111010111110111111111111100011",
8394 => "00000001111110110000000111111101",
8395 => "00000000111110010000110011111110",
8396 => "11111000111111111111010111111110",
8397 => "11110010111110011111111011011111",
8398 => "11111011000001111110000011111011",
8399 => "11011010111101111111000111101111",
8400 => "00000011111110111111010100001000",
8401 => "00000001111101110000001111111000",
8402 => "00000111111011101111110111111010",
8403 => "00010000000001100001100111111110",
8404 => "11110010000000010000011011111000",
8405 => "11111101000001111111100111101110",
8406 => "11110000111111001111001011111101",
8407 => "11011111111101101111010000000011",
8408 => "11100101111111001111101100001100",
8409 => "11111101000000001111110100000100",
8410 => "00001110111010100000010011111001",
8411 => "00000101000101111111111000000010",
8412 => "11101011000000100000000011101100",
8413 => "11111101000100100000011011101011",
8414 => "00000101111100011111000111101001",
8415 => "11100010111101110000100011111110",
8416 => "11111100000001011111101100000001",
8417 => "11111101000001000000000111111110",
8418 => "00001011111111101111101111101101",
8419 => "11111111111111111111110000000001",
8420 => "11101010111101111111110011100111",
8421 => "00000001000000110000001011100100",
8422 => "11111101111111101111010011110001",
8423 => "11101111111110101111011011110100",
8424 => "11110100000000111111101111111011",
8425 => "00000010111101010000000011111101",
8426 => "00001010111101101111101111111000",
8427 => "11111001000010111111100000000001",
8428 => "11111011111011100000000011111010",
8429 => "11111001111111100000101011101101",
8430 => "00000101111110010000000111110100",
8431 => "11110011000000000000010011111110",
8432 => "00000101000010011111010111111110",
8433 => "00000101111110000000011111111110",
8434 => "00000110111111111111111011111111",
8435 => "11111011000010110000001000000101",
8436 => "11101010111101111111110011110001",
8437 => "00000100111111010000011100000101",
8438 => "00000011000001000000011111100100",
8439 => "11111010000001001111110111111011",
8440 => "11111011111111000000011100000010",
8441 => "00001011000000011111001000000100",
8442 => "11110111111111011111100111111001",
8443 => "11110011111111110000010011110100",
8444 => "11110010111110111111001011111011",
8445 => "11111101111101111111101111111111",
8446 => "11111100111110000000000100000000",
8447 => "11111110111100011111111011111001",
8448 => "11111100111101100000000100000010",
8449 => "11111010111101111111100111101110",
8450 => "11111001111111000000100000000101",
8451 => "11100001000000001111111011111110",
8452 => "00000000000000001110111111111110",
8453 => "11111001000000010000011011111110",
8454 => "00010010111011011111000011110000",
8455 => "11110110111111110000110100000000",
8456 => "00001101111111010000010000000010",
8457 => "00000001000001110000100111100100",
8458 => "11110100000111100000000111111011",
8459 => "11100110111110010000101011110111",
8460 => "00010010111111011110100000001001",
8461 => "00000010111100111111101000000111",
8462 => "00000000000111011110011111111011",
8463 => "00000110000001111111101000000011",
8464 => "00000111000000001110011100000011",
8465 => "11110110111111011111101111100111",
8466 => "11110101000110110000010100000011",
8467 => "11101101111111101111100100001000",
8468 => "00010011111111011101100100010100",
8469 => "11110001111110111111100111111101",
8470 => "00000010000101111101111100000000",
8471 => "11101000000001110000001111111011",
8472 => "00000110000000101111011011111101",
8473 => "00000010000001000000000011100111",
8474 => "11110010000101111111110111111000",
8475 => "11110001111010010000101111111110",
8476 => "00000100111111111101111000001001",
8477 => "11110010111100111111101011000110",
8478 => "11111010000101111100110011111111",
8479 => "11010111111111111110011011001101",
8480 => "00000000111101111110111100001000",
8481 => "11111011000000001111111011011100",
8482 => "11110110000111101111100111111100",
8483 => "11101110111010110000010011111011",
8484 => "00000111111101011101101100001010",
8485 => "11110101111010111111001111010111",
8486 => "11111111000110001011100100000000",
8487 => "11010001000000111110101111010111",
8488 => "00001110111101101110110000001101",
8489 => "11110110111110011111110111101000",
8490 => "11101111000001011111001111111011",
8491 => "00000010111000110000010100000001",
8492 => "00001011111011111110101100001101",
8493 => "00000110111001101111010011001111",
8494 => "11110110000001101100010100010101",
8495 => "10101101111110111110100111100111",
8496 => "11111110111011111111000000010010",
8497 => "11110011111111011111101011110010",
8498 => "11111001111110001111010000000101",
8499 => "00001110111010100010000111110101",
8500 => "11111010111100010000011011111000",
8501 => "11110100111101001110111011011111",
8502 => "11101100000100011110011000011110",
8503 => "10110111111110001110111111111010",
8504 => "11110111111101111111110100011001",
8505 => "11110011111101111111010011111110",
8506 => "11111100110111111110101100000100",
8507 => "00010100111011000001111111111001",
8508 => "11110111111011000000110111111100",
8509 => "00010000111100111111100000000010",
8510 => "11100010111111000000001100010100",
8511 => "11001010111110011110011100000100",
8512 => "11101010111100111111100000010100",
8513 => "11111000111110001111000100001111",
8514 => "00000111110110011111100000000001",
8515 => "00001111111110000001110011111010",
8516 => "11100110111100100001010011111110",
8517 => "11111011111110011111101000001100",
8518 => "11111001111010110000000000000101",
8519 => "11100100111100101111101000001111",
8520 => "11111010111110111111101000001001",
8521 => "00000010111111101111101000001100",
8522 => "00000001111110111111100011111010",
8523 => "00010000000000110001010111110110",
8524 => "11010000111110100001100011010101",
8525 => "00001010000010001111110011111101",
8526 => "00000001111110000000101011110000",
8527 => "00000011111011101111100100001111",
8528 => "00000100111110001111110000000000",
8529 => "00000010111011001111101100010010",
8530 => "00000000111110101111000111101101",
8531 => "00001110000000010001001011110011",
8532 => "11010100111010010001000111100011",
8533 => "00000001000001110000000000010000",
8534 => "00000000111110111111011011011101",
8535 => "11111000111100101111100000010000",
8536 => "00000010111100111110110000000010",
8537 => "11111100111100101111010100010110",
8538 => "11111001111101101111101011011101",
8539 => "11111100111111010000010111110101",
8540 => "11100100110011100000000111110011",
8541 => "11111110111101001111110000000111",
8542 => "11111010111101101101101011101111",
8543 => "11011000111011011111011100000110",
8544 => "11110001111010001101101111111110",
8545 => "11111010111011111111110100000010",
8546 => "11110101000000011111100111110010",
8547 => "11101111111101000000001011110110",
8548 => "11101010111100101111010011110101",
8549 => "00000100111101101111110011111100",
8550 => "11110110111110011111101111110111",
8551 => "11110101111100111111010111110001",
8552 => "11111011111101011111110000000000",
8553 => "11110101111110011111110011110110",
8554 => "00000111111101010000001111110011",
8555 => "11011100111111101111111111111111",
8556 => "11110111000000001111100111111011",
8557 => "11111101111111101111111011111001",
8558 => "00001001000000101110111111110000",
8559 => "11100111111101100000101011111011",
8560 => "00001001111111001101001011111110",
8561 => "11111111111110011111111011101010",
8562 => "11111011000100010000000011111000",
8563 => "11100101111101011111110111111100",
8564 => "00001111111110111110010000001011",
8565 => "11111011111101001111010011111101",
8566 => "00000001000110001110011011111000",
8567 => "00000000000010101111100111111001",
8568 => "00000111111111011110111000000010",
8569 => "11111100000000000000001111101000",
8570 => "11111101000111001111110100000101",
8571 => "11101000111111111111110111111111",
8572 => "00010100000000001101111100010110",
8573 => "11110110111110000000000011110010",
8574 => "00000001000100011110101100000000",
8575 => "11110011000000110000010111111001",
8576 => "00000111111111101111110111111100",
8577 => "11111011000001100000000111011010",
8578 => "11111010000100101111110011111011",
8579 => "11101010111100011111101100000001",
8580 => "00000101111111111100010000001001",
8581 => "11111010111101000000000111011010",
8582 => "11111101000100001101111000000010",
8583 => "11101000111111011111101111100011",
8584 => "11110111000000101111110100001001",
8585 => "11111101111111011111110011001001",
8586 => "11101000000010001111011100000001",
8587 => "11101010111001011111110100000101",
8588 => "00000111111111101100111000001011",
8589 => "11110001111010101111101010111001",
8590 => "11111001000001001101011100011000",
8591 => "11100000111111101110010111000111",
8592 => "00000100111110111111100100010100",
8593 => "11111101111110010000001111101111",
8594 => "11101011000100001110111100000010",
8595 => "11111100110110000001100100000100",
8596 => "00000101111101001110011100000111",
8597 => "11110101110111111110110011001101",
8598 => "11111001000101001111001000100000",
8599 => "11100010111111001101100111001001",
8600 => "00000010111011000001000100010110",
8601 => "11110011111100101111101111110000",
8602 => "11110001111101111110110000000110",
8603 => "00001011111001110010010111110010",
8604 => "11110000111100100000010011110110",
8605 => "00100001111011001111001011101001",
8606 => "11100101000010110001011100100111",
8607 => "11101010111100011101010011101111",
8608 => "11101101111010010001001100101010",
8609 => "11110001111011111111010100000100",
8610 => "11110000110110011110110011110001",
8611 => "00001010111011110001010111101111",
8612 => "11100100111010010000100111100010",
8613 => "00100100111011101111011100000000",
8614 => "11011000111001110001010100100000",
8615 => "11101000111010011101110011111011",
8616 => "11011000111100000000001100101100",
8617 => "11110111111100111111001100000010",
8618 => "11111111110011001111000011110110",
8619 => "00001011111111100000111111110101",
8620 => "11001111111100110001010011011000",
8621 => "00011000000000110000001100010010",
8622 => "11110011110101000001101111110101",
8623 => "11110101110110111111100100001101",
8624 => "11100111111110100000100100011000",
8625 => "00000001111100011111010100001110",
8626 => "00000100111010101111100111110100",
8627 => "00000011111111100001001011110010",
8628 => "11001110111011010001011111001010",
8629 => "00000101000001001111101100010000",
8630 => "00000010111100010000011111111001",
8631 => "00000001111000111111110100001101",
8632 => "11111100111110100000000000001011",
8633 => "11110101111101001111010100001010",
8634 => "11111111111100111111110011111100",
8635 => "11101001111111011111001011110100",
8636 => "11101111111100011111101011110101",
8637 => "00001000111101001111101100000110",
8638 => "11111010111010100000010011111110",
8639 => "11111001111011110000000011111101",
8640 => "11110110000000100000000100000111",
8641 => "11111101111111011111011011110000",
8642 => "11101001111100111111001111110110",
8643 => "11010101111001111110000011110111",
8644 => "00000001110110001100110100000100",
8645 => "00000100110101001111001111111100",
8646 => "11101011111100101111110111101000",
8647 => "11111001111110111101010011011100",
8648 => "11101110111001101111111000000100",
8649 => "11110010111101011111001011010010",
8650 => "11110100111111011111010111110010",
8651 => "11110110111100101111111011110110",
8652 => "11100110111101101110111111101111",
8653 => "11111101111010111111001011111100",
8654 => "11111000111110101111110011110100",
8655 => "00000000111011011110110111100110",
8656 => "11110111111100110000000111111101",
8657 => "11110100111100001111100111101100",
8658 => "00000001111100110000001111110111",
8659 => "11010110000001011111011111111111",
8660 => "00000000111110101101110011111101",
8661 => "11111110000001100000000011111000",
8662 => "00000010111100011110010111101111",
8663 => "11011011000000010000010011110111",
8664 => "11111101111111111101010000000000",
8665 => "11111110111111111111100111011010",
8666 => "11110111000111110000000100000110",
8667 => "11100110111111011110010011111010",
8668 => "00010000000011001101100000010010",
8669 => "11110011000000000000000011110101",
8670 => "00001100000101011110010011111000",
8671 => "00000011000011000000100111110101",
8672 => "00001110000000110000000111111011",
8673 => "00000000000001011111111011100111",
8674 => "11111010000101010000001100001000",
8675 => "11100110000010111111110000000111",
8676 => "00010011000000001101100100010101",
8677 => "11100000000011110000011111110110",
8678 => "00000100000101111110011011111001",
8679 => "11111001000011010000101111111001",
8680 => "00000010000000101111101111110101",
8681 => "00000000000001100000010011100111",
8682 => "11111001000011101111110100000010",
8683 => "11011001111110111110101111111110",
8684 => "00000010000010011011000000000111",
8685 => "11100011111111100000011010111110",
8686 => "00000010000001111110001111110001",
8687 => "11111001000000101111110111010100",
8688 => "11111111111111101111010000000011",
8689 => "00000001000000010000001111000110",
8690 => "11110111000001111111111000000000",
8691 => "11110010111010111111110000001000",
8692 => "00000010111110011101100100001010",
8693 => "11100100111110000000001010111110",
8694 => "00000011000010001101001011111111",
8695 => "11100000000000101110110111010111",
8696 => "11111110111101111111101000001110",
8697 => "00000100111101110000010011100110",
8698 => "11110111000000101111111111111110",
8699 => "11111111111101000000100011111010",
8700 => "11110001111110111110010111110111",
8701 => "11111000111101001111101011010000",
8702 => "11111101000000111111010100010010",
8703 => "11110100111011001111001011010111",
8704 => "11111101111110110000000000010010",
8705 => "11111101111100001111111111110101",
8706 => "11110100111011011110111011111111",
8707 => "00001011111110100001011011101111",
8708 => "11101000000000000000011011101001",
8709 => "00100100111110111110110011101110",
8710 => "11101100111101000010011000011100",
8711 => "00000100111010101110110011111111",
8712 => "11101010111100110001011000010010",
8713 => "11111000111100101111001000000101",
8714 => "00000010110111101110111000000001",
8715 => "00001110000001100000001011110011",
8716 => "11011001111110110001100011011010",
8717 => "00101101000001101111110011111111",
8718 => "11101000110100110010101000000001",
8719 => "00001110111001101111100000001011",
8720 => "11101110111111100001111100010011",
8721 => "11111101111101011111000100001010",
8722 => "00000001110110101111110000001000",
8723 => "00000100000011000000000111110111",
8724 => "11100010111011100001100011100011",
8725 => "00011001000001010000000000000111",
8726 => "11110010110110000010000011110011",
8727 => "00000010111010110000101100001100",
8728 => "11101101000010010001011100000111",
8729 => "11111110000000111111010000001000",
8730 => "00000001111101100000010000001001",
8731 => "11110110000010011110011011111110",
8732 => "11101001000000111111111111101000",
8733 => "00001000000001101111111011111001",
8734 => "11111010111001110001110000000001",
8735 => "00010010111101110000011100001111",
8736 => "11111011000000010001001000000110",
8737 => "11111101000011111111110000000010",
8738 => "00000011111111100000001100010001",
8739 => "11100110000100011101000000000001",
8740 => "11110010000010011101101011111111",
8741 => "00000000000100010000110111111101",
8742 => "11111101111010110000100011100011",
8743 => "00001100000000000000011111110001",
8744 => "00000011000010000000100011111101",
8745 => "00000111000010100000001011101110",
8746 => "11111000000011011111010000000011",
8747 => "11110000111010001110100111111100",
8748 => "11111111111111111101111111111001",
8749 => "00000001111110111111100111111001",
8750 => "11110001000010110000011111100111",
8751 => "00001000111110111110110011011111",
8752 => "11110101111010100000111100000001",
8753 => "00000000111101111111011111100011",
8754 => "11110010000000011111100111110011",
8755 => "11100111111011111111110011110110",
8756 => "11011011111101101110010111100110",
8757 => "00000010111100101111001011111001",
8758 => "11111100111110100000000111111011",
8759 => "00000000111001111111011011100111",
8760 => "11111111111011000000001111111111",
8761 => "11110010111011111111000111101010",
8762 => "00001011111011100000001111111001",
8763 => "11100100000001001110111111111100",
8764 => "00000111111111001111001000000000",
8765 => "00000001000001010000001000000000",
8766 => "11111010111101001110110111110010",
8767 => "11011011000010000000001000000011",
8768 => "11101110000000101101110100000100",
8769 => "00000100000001101111110011110011",
8770 => "00000111001010010000100011111101",
8771 => "11101000000001011101101000000000",
8772 => "00000101000010001110111100001010",
8773 => "11111000000000111111110011110001",
8774 => "00010001001001011101100011111100",
8775 => "00001111000001000001011111111011",
8776 => "00001010000000101110111111110111",
8777 => "11111101000001010000011011110110",
8778 => "00000001000101000000010000000100",
8779 => "11100011000000111110000100001100",
8780 => "00001101000001011101100000010010",
8781 => "11100100000001100000010111101101",
8782 => "00000110000100111101100011110111",
8783 => "11110011000010110000010111110111",
8784 => "00001000000001101111111111111010",
8785 => "00000010000100110000010011100000",
8786 => "00000101000100000000101011111101",
8787 => "11010000000010111101010111111111",
8788 => "00001110000000101011100000001100",
8789 => "11011101000010110000101011000110",
8790 => "00001101000001011101000111101011",
8791 => "11100010000001110000111111100101",
8792 => "00000000000011011110011111110001",
8793 => "00001001000001110000101011000101",
8794 => "00000000000010000000101100000010",
8795 => "11100101111111111110010011111110",
8796 => "00000100000000111100100000000011",
8797 => "11101100111110100000000010111100",
8798 => "00010000111110111110000111111010",
8799 => "11110110000000010000010011001011",
8800 => "00001101000001111111110111110011",
8801 => "00000011111111010000011111011000",
8802 => "11101001000010111111001100001100",
8803 => "00000011111100000000100000000100",
8804 => "00000000000000001110111011111001",
8805 => "11111000111011111111010111010100",
8806 => "11110110000010100000011100101001",
8807 => "11111001111111011110010011101000",
8808 => "00001011111101100001000111111011",
8809 => "11111101111110010000001011110000",
8810 => "00000111111101111111010100010001",
8811 => "00010001000000000001010011110110",
8812 => "00001110000000100001010100001011",
8813 => "00001001000001011111010100000000",
8814 => "11111011000000010010100000101110",
8815 => "00011010000000100000010000001111",
8816 => "11111110000000110010000000000100",
8817 => "00000011000001011111001100010101",
8818 => "00001101111100010000011100000101",
8819 => "11110110000011111101100111111000",
8820 => "11111000000010000000011111110010",
8821 => "00100100000010010000001011111011",
8822 => "11111111110111000001111100001101",
8823 => "00011010111111010000110100001101",
8824 => "11101111000011100001100111111110",
8825 => "00000001000011001111101100000000",
8826 => "11111110111101101111111100000011",
8827 => "11101010000000111101000000000010",
8828 => "11110011000010111111000111111010",
8829 => "00000101111111001111111111111101",
8830 => "00000100111000000001010111110110",
8831 => "00001111111111000000001000000000",
8832 => "11111101000000000000110011111100",
8833 => "11111011000000000000001011101100",
8834 => "11111111000000100000010100001001",
8835 => "11110110000011001110010000000100",
8836 => "11111111000100011111100111111110",
8837 => "00000011000100010000101100000101",
8838 => "00001000111011100000010011100101",
8839 => "00000110000000010000010111111101",
8840 => "11111111000000010001001111111011",
8841 => "00001011000001010000001111111001",
8842 => "00000101000010010000010000001001",
8843 => "11111011111111101111110100001010",
8844 => "00000101000001111111100000000111",
8845 => "00000101000000100000011100001011",
8846 => "00000111000010011111110111011101",
8847 => "00001000000000101111111100001011",
8848 => "00001000000000000000001011111010",
8849 => "00000111000010100000111000000001",
8850 => "11111110000011111111111000000010",
8851 => "00000101111110010000000011111101",
8852 => "11101001111100001110111111101110",
8853 => "00000101111111010000001111111111",
8854 => "11111100000010010000000111111010",
8855 => "00000001111111101111000111110000",
8856 => "00010000111110101111111000000000",
8857 => "00000010111110001111111111110101",
8858 => "11110100111111011111001111111001",
8859 => "11101011111110010000010011110100",
8860 => "11011110111101001110011111101010",
8861 => "00000000111110001111100111111001",
8862 => "11111000111101110000000000000001",
8863 => "00000011111000111111010111101100",
8864 => "11111110111101110000010100000010",
8865 => "11110110111110001111011011100111",
8866 => "00000011111101001111010111111110",
8867 => "11101010111101001110110011111111",
8868 => "00010000111111011110111000001000",
8869 => "00000000000001110000001000000001",
8870 => "11101000111010111111011111111010",
8871 => "11100001000001111110110000000110",
8872 => "11101000111110001110111000000100",
8873 => "11111111000010101111010011110001",
8874 => "00000010001000110000010100000001",
8875 => "11101100000011001101011100000100",
8876 => "00010000000001001111100100010100",
8877 => "11111101000001001111110100000110",
8878 => "00001101000100111101001111110100",
8879 => "00001001000011000000111000001010",
8880 => "00010000000000001111011011111111",
8881 => "00000111000000100000000011111010",
8882 => "00000000000101010000010000001101",
8883 => "11011001000011001110010100000101",
8884 => "00001101000000111101111000010000",
8885 => "11010100000010010000100111110101",
8886 => "00001110000100111110110111110100",
8887 => "11111101000011100000100111111010",
8888 => "00001010000010010000000011110111",
8889 => "00001101000010010000011111100100",
8890 => "00000100000011010000011000000111",
8891 => "11011011111110111100101100001011",
8892 => "00011110000010001101011000011001",
8893 => "11100100000000100000100011100101",
8894 => "00010000000000101100111011011101",
8895 => "11100100000011100000100111101100",
8896 => "00000011000010111110111011100000",
8897 => "00001001000100000000011111011100",
8898 => "00000011000101100000101111111000",
8899 => "11110001000010001110111000000000",
8900 => "00001010000000011110010000010010",
8901 => "11100110000010100000011111011010",
8902 => "00010011111111111101100111101001",
8903 => "11110111000000110001101111101101",
8904 => "00010101000010011101111011011111",
8905 => "00001000000001110000011011101011",
8906 => "11111111001000101111111100000001",
8907 => "11111001000001000000001111111111",
8908 => "00000100000011001111011000000000",
8909 => "11110101000000110000000111110111",
8910 => "00001001000101000000101000010110",
8911 => "00100101111111111111110011111010",
8912 => "00010010111111000000011111101000",
8913 => "00000110111011100000000111111100",
8914 => "00000100000100001111111000001010",
8915 => "00000000000010011111100111111110",
8916 => "00001001000011110000010100001110",
8917 => "00000111000000110000000000010000",
8918 => "00000000111101110001111000001110",
8919 => "00100101000001110000010100001011",
8920 => "00001010111111100001111011100000",
8921 => "00000011111111110000010000000101",
8922 => "00000010000010111111111100000011",
8923 => "00000011000100101111100100000000",
8924 => "00000000000010100000011011111101",
8925 => "00011011000011001111111111111111",
8926 => "11111111111110100001111011111111",
8927 => "00010010111111110000101000000101",
8928 => "00000010000010110001011011110010",
8929 => "00000011000000100000001000001000",
8930 => "00010010000011100000011000000101",
8931 => "00001100000011000000100111111110",
8932 => "11111101111111100001000000000011",
8933 => "00000101000011000000001111111101",
8934 => "00000111000001110000110100000100",
8935 => "00000111000000100000101100001010",
8936 => "00001110000010110001100011110011",
8937 => "00000010000001110000101000001001",
8938 => "00001001000010010000010111111011",
8939 => "00001101000011110000101011111110",
8940 => "00001111000001010000010100001010",
8941 => "11111110000010110000100100000001",
8942 => "00001100000000101111000000000010",
8943 => "11110110000000110000111000000100",
8944 => "00000011000011010000100011111010",
8945 => "00000010000001110001000000000011",
8946 => "00001011000000010000101111101101",
8947 => "00000001000010010000001011111110",
8948 => "11111101000001000000011011111001",
8949 => "00000000000010100000100011111011",
8950 => "11111111000000001111100100001010",
8951 => "11111001111111100000000100000100",
8952 => "00000000000001111111110111111011",
8953 => "00001001000001010000010000000010",
8954 => "11111111000001001111111111110000",
8955 => "11111111000000001111101111111000",
8956 => "11100000000000011111010011100110",
8957 => "00000111111101100000000011111101",
8958 => "00001110111111100000011011110011",
8959 => "11111100111101011111101111110011",
8960 => "00010101111110101111110011111101",
8961 => "00000101111110010000100011110001",
8962 => "11110110111111011111010111111011",
8963 => "11101000111110010000001011110110",
8964 => "11101010111101101110101111110110",
8965 => "11111100111101011111010111111110",
8966 => "11110101111101110000001111111110",
8967 => "00000010111101111111100111110001",
8968 => "11111111111110010000010000000010",
8969 => "11110110111111001111100011101010",
8970 => "11110000111111011111010000000011",
8971 => "11111010111010101111000111111011",
8972 => "00000101111110011111100000001110",
8973 => "11111101111110011111011100001011",
8974 => "11110001000000001111010111110101",
8975 => "11101000000010101111001000001010",
8976 => "11111010111110010000010100000110",
8977 => "11110101000000011111111011101110",
8978 => "11111110000010101111111011111101",
8979 => "11110101111111111110101011111001",
8980 => "00001101111110111111100100001111",
8981 => "00000100111110111111110000010001",
8982 => "00000011111111111101010011100100",
8983 => "11110000000001110000011100000111",
8984 => "00000001000000001110011100000101",
8985 => "00000011111111110000000011110101",
8986 => "00001000000100000000110100000001",
8987 => "11100111000011011101110000000011",
8988 => "00010001000010001111010100010000",
8989 => "11101101000010000000001100000110",
8990 => "00001100000010111110001011011011",
8991 => "11111100000011110000111100000110",
8992 => "00000111000001011111011111101000",
8993 => "00001000000010000000101111110010",
8994 => "00010000000111010000011111111010",
8995 => "11100111000001101100110100001101",
8996 => "00001110000010011110101000010001",
8997 => "11100101000010110000101000000000",
8998 => "00001110000101011101101111010100",
8999 => "11110101000010000001000100000100",
9000 => "00010011000010111110011111010100",
9001 => "00000101000010110000100011110000",
9002 => "00000011000100110000010100000011",
9003 => "11101000000000111101010100001001",
9004 => "00010010000001001110101000010110",
9005 => "11001101000000010000111100000000",
9006 => "00010011000010001110000111101001",
9007 => "11111110000100110000110111111101",
9008 => "00001100000011001110110111010011",
9009 => "00000101000010110000101011110000",
9010 => "00000011000101110000100000000100",
9011 => "11110001000010111110010000000010",
9012 => "00000000000001101110010111111010",
9013 => "11111101000010110000101011110010",
9014 => "00000001111110101111000011101010",
9015 => "00000001111110101111101111101000",
9016 => "00001111000000011111111111110000",
9017 => "00010000000000110000000111110000",
9018 => "11111111000110100000011000000000",
9019 => "00000000000000111111101111111111",
9020 => "00000110000010111111011100000101",
9021 => "00000000000000100000010100001010",
9022 => "00000101000001111111101111101100",
9023 => "00010101000000111111111100000000",
9024 => "00001011000010010000110011011011",
9025 => "00000010000001010000100011111110",
9026 => "00000111000100000000100011111001",
9027 => "00001011000000000001000100000101",
9028 => "00000010000000110000111000000011",
9029 => "00000000000001100000010000001000",
9030 => "00000101000100100000011100000110",
9031 => "00001110000001000000011000000110",
9032 => "00000001000100000000001111101100",
9033 => "00001010000001100000011100000111",
9034 => "00000101000010001111110111111001",
9035 => "00001001111111100000110000000011",
9036 => "11111111000001110001000111111001",
9037 => "11101111000001011111111000000010",
9038 => "00001001000011110000001000000100",
9039 => "00001001000001000000001000000101",
9040 => "00000111000001100001010011110010",
9041 => "00000000111110101111111000001011",
9042 => "00000100111111110000010111111011",
9043 => "00000011000001100000000011111111",
9044 => "11111001111111111111101100000011",
9045 => "00001110111110010000000100000000",
9046 => "00000000111111111111100011101111",
9047 => "11101100111111000000011111111010",
9048 => "11111111000001110000011011111001",
9049 => "11111110111111001111110111111101",
9050 => "00000100111110000000000111110110",
9051 => "00001001000001000000000000000001",
9052 => "00000010111110010000010100001000",
9053 => "00000000000010000000011100000001",
9054 => "00000001111111011111101100000001",
9055 => "11110101111111111111110000010001",
9056 => "00000010000000110000000100000001",
9057 => "00000110000000010000011000001100",
9058 => "00001010111111010000001011110101",
9059 => "00001000000011000000001011111000",
9060 => "11101110111101100000001011110111",
9061 => "11111001000001100000010011110110",
9062 => "00000101111111101110101011111111",
9063 => "11110101111100100000011100000111",
9064 => "00001100000001011110010011111100",
9065 => "00001011111101111111111000000110",
9066 => "11111001111111001111010011111001",
9067 => "11101011111111000000000111111000",
9068 => "11110001111101001110100111111010",
9069 => "00000000111101001111101000000010",
9070 => "11111011111110100000001011111101",
9071 => "11111111111101011111110011110001",
9072 => "11111011111110000000001100000001",
9073 => "11111011111110011111100111110010",
9074 => "11110010000000011111100111111000",
9075 => "00001001111110000000011011111001",
9076 => "00000000111110000000010100000010",
9077 => "11111101111111101111101000000111",
9078 => "11111001111111011111111011101010",
9079 => "11110100111111001111100000000000",
9080 => "11111010111101100000011100000001",
9081 => "11111001111110101111100000001010",
9082 => "00000010111100101111110111110110",
9083 => "11111110000001001110111111111100",
9084 => "11111110111111011111101000000001",
9085 => "11111101000010001111111000000111",
9086 => "11111100111010111110100111011011",
9087 => "11101101111101111111110100000011",
9088 => "11110001000000111111110111111110",
9089 => "00000011111111111111100011111110",
9090 => "00001011000100110000011011110101",
9091 => "11110101000000101110101100000011",
9092 => "00000100111111100000000000000011",
9093 => "00001001000001101111111100001111",
9094 => "00000100111100111110010111001100",
9095 => "00000000000001110000101100001101",
9096 => "00000110000001101110111011111110",
9097 => "11111101000001010000100000000011",
9098 => "00001000000101110000011111111011",
9099 => "11101111000001111110001000000110",
9100 => "00000111000000111111110100001010",
9101 => "00001000000010010000110000010010",
9102 => "00001001000011101110101011001111",
9103 => "11111010000001110000110100001001",
9104 => "00001001000010111111100011100011",
9105 => "00001101000011010000001100000000",
9106 => "00010000000010110000110111110010",
9107 => "11111100000101101101111000000110",
9108 => "11110101000000110000100111111011",
9109 => "00001101000010110000011100011100",
9110 => "00010000111111011110111111010011",
9111 => "11111111000000110001110100001010",
9112 => "00001000000011011111001111001111",
9113 => "00001000000010110000100000001001",
9114 => "00010001000001000000110011110110",
9115 => "00000010000110001110110100000001",
9116 => "11100010111111000000000011100010",
9117 => "11111100000001110000100000001101",
9118 => "00000111111000101111010111110000",
9119 => "00001000111101010001011000001000",
9120 => "00000011000100001111111111100001",
9121 => "00001010000001110000010100000111",
9122 => "00001000000011100000110011111011",
9123 => "00001110000010100000101000000000",
9124 => "11101011000000100000101011101000",
9125 => "11101100000010110000010011111010",
9126 => "00000001000011101111011111111010",
9127 => "00000100111110010000000111111101",
9128 => "00000101000010001111111011011100",
9129 => "00001000111111010000100100000100",
9130 => "00000011000001000000100111111101",
9131 => "00010100000001100001010100001000",
9132 => "11110110000000110000111111110101",
9133 => "11100100000011001111111011101001",
9134 => "11111111000100001111000100010001",
9135 => "00000001111111000000010100000101",
9136 => "00000000000000000000010111110110",
9137 => "00000110000000100000001000001011",
9138 => "11111111000000100000010000000001",
9139 => "11111111111111110000010011110111",
9140 => "00000100000001100000001011111111",
9141 => "11111101000000100000000011110010",
9142 => "11111100000001010000001000011011",
9143 => "00000010111111001111111100000101",
9144 => "00001001111111110000000111111010",
9145 => "00000100000001010000001100000101",
9146 => "00000010111101100000010011111100",
9147 => "11111110111111101111110100000010",
9148 => "11100110111101111111111011101110",
9149 => "11110110111111110000010011101100",
9150 => "00000001111111111111100011110110",
9151 => "11111000111101001111101011111100",
9152 => "00000100000001001111110100000001",
9153 => "00000100000000010000010000000000",
9154 => "00000111111110011111101111111100",
9155 => "00000000000000110000011111111000",
9156 => "11110010000000110000010111110001",
9157 => "11111110111111000000001011111000",
9158 => "11111001111111010000011000001101",
9159 => "11111010111110011111110000000011",
9160 => "11111110111111011111111011111111",
9161 => "00000010111110101111110000000011",
9162 => "00000000111110000000000011111001",
9163 => "00000011111110110000001011111110",
9164 => "00000010111101110000010111111101",
9165 => "11111110111110111111111011111111",
9166 => "11111110111111111111010011111000",
9167 => "11110100111110100000010100000011",
9168 => "00000000000000011110101111111111",
9169 => "11111100111111001111110100000101",
9170 => "11111101111110101111101111111101",
9171 => "11110010111110110000001111110111",
9172 => "11110101111110111111000011111100",
9173 => "11111110111101111111110011111110",
9174 => "11111011111101101111111000000000",
9175 => "00000011111110101111100111110111",
9176 => "11111011111110010000000011111101",
9177 => "11111001111110011111011011110111",
9178 => "11110111111111011111101011110100",
9179 => "11111101111100110000110111110111",
9180 => "11011101111100010000000011101010",
9181 => "11111101111100011111011111111011",
9182 => "11111000111101110000001011111011",
9183 => "00000001111011101111011011110110",
9184 => "11110100111110001110111011111111",
9185 => "11110111111101101111001111110111",
9186 => "11110111111110111111001011110011",
9187 => "00000011111010101111111011110110",
9188 => "11111000111011100000011011111011",
9189 => "11111111111100001111010000001110",
9190 => "11101101000000001111110111110110",
9191 => "11110000111110001110011100000101",
9192 => "11110001111010011110100000000101",
9193 => "11101100111111011111110100000100",
9194 => "00001000111010110000101011110111",
9195 => "11111110000000001111101011111101",
9196 => "00000110111110110000000000000001",
9197 => "11111110000000111111101100001010",
9198 => "00001011111101001101111111100111",
9199 => "11101000000010010000101000000011",
9200 => "00001001111111111110100100000000",
9201 => "11111000000000000000011111111100",
9202 => "00001001000010000000110011101110",
9203 => "00000100000001011111100011111101",
9204 => "11111100111101010000010011111100",
9205 => "11111111000010010000111100001110",
9206 => "00001001111111011101100111010101",
9207 => "11110100000001010000101000000100",
9208 => "00001100000011101110011111111001",
9209 => "00000000000001000000001000000010",
9210 => "00001000000001100000010111110010",
9211 => "00001000000010001111011000000110",
9212 => "11110101111100110000100111110001",
9213 => "00010011000001000000100100010010",
9214 => "00000111111011011111111011100011",
9215 => "00001000000001000000111000001100",
9216 => "11110101000011111111100011110111",
9217 => "00000100000000000000000100010000",
9218 => "00001000111111010000000011111001",
9219 => "00000101000111110000100000000100",
9220 => "11010110111111100001010111010101",
9221 => "00100010000011010000100000000111",
9222 => "00000001111101010000011011010100",
9223 => "00000110111110000000110100010011",
9224 => "00000101000000010000101011010101",
9225 => "00001000000000110000001100001111",
9226 => "00000001000001100000010011111100",
9227 => "00010010000100100001000011111101",
9228 => "11010110000000000001000011011000",
9229 => "00001010000000110000000100000110",
9230 => "11111001000100000000101000010111",
9231 => "00010010111011111111101100001111",
9232 => "00000001111111010000001011111001",
9233 => "00000000111111010000000100010010",
9234 => "11111111111111000000000100001111",
9235 => "00001101000001110000101100000000",
9236 => "11111010000010100000100111110111",
9237 => "11101101000010101111101011111000",
9238 => "11111010000000010001001000011001",
9239 => "00000100111110111111111000001000",
9240 => "00000001111111000001001000000010",
9241 => "00000000000001110000010000001111",
9242 => "11111110111110101111011000000011",
9243 => "00000010111111110000010000000011",
9244 => "11110010000001111111110011111110",
9245 => "11101111000000001111101011100101",
9246 => "11110111000000010000001000001010",
9247 => "11111011111111011111101111111010",
9248 => "11111001111111000000101111111110",
9249 => "11111011111111000000000011111010",
9250 => "00000010000000011111101011111001",
9251 => "00000001111110110000000111111111",
9252 => "11110001111110001111110111110100",
9253 => "11111011000011011111101111100110",
9254 => "00000101000000111110001100000011",
9255 => "11111000111100001111010111111010",
9256 => "11111111000001001111001000000110",
9257 => "11111101111111110000000011111011",
9258 => "11111001111101101111011011101111",
9259 => "11111001111011110000000011110110",
9260 => "11011001111011011111100111101110",
9261 => "11111111111100001111110011110111",
9262 => "11110010111111111111010100000100",
9263 => "11110000111100111110111011110011",
9264 => "11101101111011001101101000000010",
9265 => "11110001111100111111111011110100",
9266 => "00000001111010011111011011110110",
9267 => "00000000000000001111111111111000",
9268 => "00000010111100100000011100000001",
9269 => "00000000111111101111110000000011",
9270 => "11110100111011111111000111111111",
9271 => "11010100111111000000001000000101",
9272 => "11110100000000111110101011111110",
9273 => "11110100111110001111010100000101",
9274 => "11111111000000000000000111111111",
9275 => "00000000000000110000000011111011",
9276 => "11111100111111100000000100000000",
9277 => "00000011111111111111110111111111",
9278 => "11111100111110110000001111111111",
9279 => "00000010111110100000000100000001",
9280 => "00000001000000010000011111111101",
9281 => "00000000000000011111111111111101",
9282 => "11111001111111111111010011110011",
9283 => "11010010111110001111011111110010",
9284 => "11010111111101011101010011101101",
9285 => "00000000111100111111011111110010",
9286 => "11110111111110101111110100000011",
9287 => "00000001111011111111100011100011",
9288 => "11110100111110011111110000000000",
9289 => "11110110111101111111100011100000",
9290 => "11101110111111001111000111110101",
9291 => "11011011111001001110101011101110",
9292 => "11110001111100011110001011110101",
9293 => "11111100111100101111001011110100",
9294 => "11101101111000110000000111111101",
9295 => "00000011111101101110010111011110",
9296 => "11101111111100001111111000000101",
9297 => "11110000111011001110111111010111",
9298 => "11111010111100011111100011101110",
9299 => "11111100111110111111101011111011",
9300 => "11111110111101000000000000000101",
9301 => "00001110111101111111101100001001",
9302 => "11110111111011001111111111111010",
9303 => "11111111000001111111101011111010",
9304 => "11111000111100011111100000000100",
9305 => "11111101111111111111100011111001",
9306 => "00001010111111110000100111110010",
9307 => "11111110000001000000001111111101",
9308 => "11101001000000010000100111110100",
9309 => "00000111000001101111110000001100",
9310 => "11111001000011110000010000000001",
9311 => "00000100111100010000000000000011",
9312 => "00000010111110001101011000001001",
9313 => "11111111111110111111100011111101",
9314 => "00001110111010110001000011110011",
9315 => "00000001000000110000000111111100",
9316 => "11011010111110110000100111101111",
9317 => "00001010000001100000000100001101",
9318 => "00000101111101011111110111110111",
9319 => "11101111111100100000001100001011",
9320 => "11110011000000101100100011111101",
9321 => "11111110000000110000010011111111",
9322 => "00000100110111101111111111101111",
9323 => "00000001000010110000001111110110",
9324 => "11001101111110000000001111011001",
9325 => "00000001000001000000000000000101",
9326 => "11111000111100011110010111101010",
9327 => "11001111111010100000011000000011",
9328 => "11110110000000111101100011111011",
9329 => "00000010111111000000001000000001",
9330 => "00000001111011011111101111101111",
9331 => "11111010000001000000001011111100",
9332 => "10110001111110001111111111001010",
9333 => "11111010000001100000011011111110",
9334 => "11111010111110011110110111111100",
9335 => "11100110110111100000100111111110",
9336 => "11111100000000101111010000001011",
9337 => "00000010111110001111110111111101",
9338 => "11111101111101011111101011111001",
9339 => "11110111000000011111111100000000",
9340 => "11001100111011110000001011011010",
9341 => "00000000111110110000000011110110",
9342 => "11111001111111001111100111110100",
9343 => "11100010111011001111101111111110",
9344 => "11111001000000011111001011111001",
9345 => "11111100111100101111111111111001",
9346 => "11111101111101011111111111110100",
9347 => "11111110111111111111111000000010",
9348 => "11010100111111001111111011011100",
9349 => "11111001111111100000000111111111",
9350 => "11111010000000001111011111111100",
9351 => "11011111111010101111100100000000",
9352 => "11111011111101111110010011111100",
9353 => "11111100111110000000001011111110",
9354 => "11111111000000111111001111101111",
9355 => "11110111111101011111110111110101",
9356 => "11001000111010111111001011100010",
9357 => "11111110111101000000000011101100",
9358 => "11110100000000111111101100001000",
9359 => "11111011110110101111101111110010",
9360 => "11111001111110001110110011111111",
9361 => "11111011111010101111101111101110",
9362 => "11101011111001001110101011111000",
9363 => "11011100111001011110010011101011",
9364 => "11100010111011001110000111101110",
9365 => "11111111111001001111010111101110",
9366 => "11101110111010001111111011110011",
9367 => "11101010111001111110101011100110",
9368 => "11110001111011001110111011111111",
9369 => "11110000111011001111011011100110",
9370 => "11101010111000001110101100000010",
9371 => "11011100111011001110111111110111",
9372 => "11111110111100001101111000000010",
9373 => "11111111111001001111001100000011",
9374 => "11101011110101100000001111110010",
9375 => "11101101111111011110100011100001",
9376 => "11101111111001000000011100000001",
9377 => "11110101111100101111010011011111",
9378 => "11111100111110111111111000000100",
9379 => "00000000111111010000000000000010",
9380 => "11111100111111010000010000000010",
9381 => "11111111111111110000000100000010",
9382 => "00000001111111011111111100000101",
9383 => "11111111000001000000001000000001",
9384 => "00000100111111010000010000000101",
9385 => "00000011000000101111110100000001",
9386 => "11111000000000001111100011111111",
9387 => "11111100111111101111111100000000",
9388 => "11111010111110001111101000000000",
9389 => "00000100111111101111101011111110",
9390 => "11111111111110010000010011111111",
9391 => "00000101111111101111100111111001",
9392 => "11111101111111110000100000000000",
9393 => "11111111111111101111101100000000",
9394 => "11110101000000001111100011111101",
9395 => "11100110111110011111110111111000",
9396 => "11100001111110001110001011110101",
9397 => "00000001111101001111011111110101",
9398 => "11110110111100110000001100000110",
9399 => "11111110111110101111100011100111",
9400 => "11111101111101111111111000000011",
9401 => "11111000111110101111010111100011",
9402 => "11110000111110011110110111111000",
9403 => "11010011111110011110111011110110",
9404 => "11010100111110101100101011101000",
9405 => "11111110111101101111100111101110",
9406 => "11110100111000100000001000000101",
9407 => "00000100111101111110100111011100",
9408 => "11110111111010110000000000000000",
9409 => "11111100111101111111010011010101",
9410 => "11110001111000001111010011110110",
9411 => "11010000111011011101101111110010",
9412 => "11101011111110001100010011110101",
9413 => "00000001111011111111011011101100",
9414 => "11110001110110000000010011110111",
9415 => "11111101111011011110001011001010",
9416 => "11110010111010011111100100000101",
9417 => "11110110111101111111100010111100",
9418 => "11111000110010100000000011111001",
9419 => "11110110111011111111001111111011",
9420 => "11101100111100111111000011111110",
9421 => "11111111111011001111100000000001",
9422 => "11110010110111000000010111110010",
9423 => "00000010111011011110010011111001",
9424 => "11110010111000100000000111111111",
9425 => "11111000111100111111100111110011",
9426 => "11111100111001100000000111111100",
9427 => "00000000111011100000000111111010",
9428 => "11111000111101001111111100000011",
9429 => "00000001111101101111110000000111",
9430 => "11111110111100110000000111111001",
9431 => "11110111111010011111101000000011",
9432 => "11110011111110001111111100000000",
9433 => "11111000111101011111100100000010",
9434 => "00000011111010010000100111111010",
9435 => "00001001111100010000110111111010",
9436 => "11100001111100110000110000000000",
9437 => "11111111111110011111110000010010",
9438 => "11111000000001000000010111101110",
9439 => "11101111111100000000011100001100",
9440 => "11111001111111011111110000000011",
9441 => "11110110111111001111111100001100",
9442 => "00001011000010000001000111110110",
9443 => "00001000111111110000101111111011",
9444 => "11011001111101010000011111101111",
9445 => "00000000111110011111111100001001",
9446 => "00000110000011110000000000000111",
9447 => "11110011111101000001001100001101",
9448 => "11111111000011010000011000000001",
9449 => "11111001000010010000010000001110",
9450 => "11111101000000110000001011111100",
9451 => "11111001111110000000010111111001",
9452 => "11101011111110001111011011110110",
9453 => "00000001111101111111010111111011",
9454 => "11110100000000110000001100000001",
9455 => "11110111111101111111111111111110",
9456 => "11110100111110100000000100000011",
9457 => "11111000000000001111101111111010",
9458 => "11101101111110111110111011111001",
9459 => "11101001111101111111011011111000",
9460 => "11111011111111001110010111111000",
9461 => "00000001111101011111101011111100",
9462 => "11101111111011100000010100000010",
9463 => "11111010111110111110100011101000",
9464 => "11110010111010010000010000000010",
9465 => "11111000111011101111011011100000",
9466 => "11110001111011011111001100000010",
9467 => "11101101111101101111100011111111",
9468 => "11111101000000001110101000000010",
9469 => "00000011111111001111101000000000",
9470 => "11111011111010101111111011111001",
9471 => "11111111000000001111000111110001",
9472 => "11111100111011110000010100000100",
9473 => "11111100111110101111100011101000",
9474 => "00000000111111101111101100000000",
9475 => "00000000111111001111111000000011",
9476 => "11111101000000011111110011111111",
9477 => "11111111000000110000000011111111",
9478 => "11111110111111000000001000000110",
9479 => "00000001000000111111110111111111",
9480 => "00000011111111100000101011111111",
9481 => "00000001000000011111101000000000",
9482 => "00000000000000000000000000000000",
9483 => "00000000000000000000000000000000",
9484 => "00000000000000000000000000000000",
9485 => "11111100000000000000001011111101",
9486 => "11111111000000110000001000000000",
9487 => "00000010111111010000010000000001",
9488 => "00000100000001000000001000000100",
9489 => "00000010000000010000001000000000",
9490 => "00000100000000110000000100000110",
9491 => "11111100111111110001100100000110",
9492 => "00000010111111010000001000000011",
9493 => "00000011000001010000001000000010",
9494 => "11111101000001001111111011111101",
9495 => "11111101000000010000001000000100",
9496 => "00000100111111110000000011111110",
9497 => "00000010000001010000001011111111",
9498 => "11111110111111010000000000000010",
9499 => "11111010111111100001101100001000",
9500 => "11111100111111101111110111111101",
9501 => "11111010111110101111101011111010",
9502 => "11111010000000111111111011111101",
9503 => "11101100111110000000001111111100",
9504 => "00000110111110111111110011111111",
9505 => "11111111000001011111111111111001",
9506 => "11111001111110101111000100000101",
9507 => "11111011111111110001010100001000",
9508 => "11111001111111011111101100000011",
9509 => "11111000111100011111101111101110",
9510 => "11111000111111001111111011111011",
9511 => "11100011111101010000011011110011",
9512 => "00000010111100011111100111111111",
9513 => "11101101111110111111011111110100",
9514 => "11101010111101011110010100000000",
9515 => "11110111111100101110101000000110",
9516 => "11110101111101111111101011111110",
9517 => "11110100111010111110111011101011",
9518 => "11110001111110010000000011110101",
9519 => "11011100111101101111110111110001",
9520 => "00001000111100001111010000000011",
9521 => "11101110111011101110111111110010",
9522 => "11011110111101001110111111111100",
9523 => "11101110111011111110011000000100",
9524 => "11111010111100111111010011110011",
9525 => "11110011110111111110111111100111",
9526 => "11110110111100111111111111110111",
9527 => "11011110111100011111110011101111",
9528 => "00000101111011101111100111111110",
9529 => "11101101111010001111000011101100",
9530 => "11010100111101011110101000000001",
9531 => "11101101111011011101101100001001",
9532 => "11110011111100111111000111111011",
9533 => "11110001110110101111000111101100",
9534 => "11111000111110001111111011110100",
9535 => "11011101111100111111111011110110",
9536 => "00001000111100011111100011111110",
9537 => "11101100111000001110101011110001",
9538 => "11010000111110101110100011111101",
9539 => "11101111111011101101101100001000",
9540 => "11110100111011101111000111111000",
9541 => "11110010111000011111011011101010",
9542 => "11110111111100101111111111111011",
9543 => "11100000111100111111111011110000",
9544 => "00000101111100011111010000000101",
9545 => "11101011111010001111000011111000",
9546 => "11010001111100101110101000000010",
9547 => "11110001111100101101111000001000",
9548 => "11111100111101101110110011110110",
9549 => "11110110110111101111101011110111",
9550 => "11110110111100000000000111110110",
9551 => "11101101111101111111111111111011",
9552 => "00000011111011001111101000000101",
9553 => "11110100111000101111011011110110",
9554 => "11010110111101101110101100000100",
9555 => "11101110111101101110001000000101",
9556 => "11111010111110111111001011111011",
9557 => "11110110111000111111100011110100",
9558 => "11111111000000100000001111110111",
9559 => "11110111111110011111111111111100",
9560 => "00001000111110001111111000000011",
9561 => "11110001111010001111111011111110",
9562 => "11100111111110111111010000000110",
9563 => "11111010111110101111010000000100",
9564 => "11111011111110111111100000000011",
9565 => "11111110111100011111111011111010",
9566 => "11111011000000001111110111110111",
9567 => "11111110111111110000000000000001",
9568 => "00000001111111011111101111111110",
9569 => "11111100111101010000000111111110",
9570 => "11111001111111011111011100000011",
9571 => "11111100111110100000101100000111",
9572 => "11111000111111011111100100000010",
9573 => "11111111111111100000000111111101",
9574 => "11111110000000111111110100000011",
9575 => "00000000111111000000000100000100",
9576 => "00001001000000011111101100000010",
9577 => "00000000111110100000010011111111",
9578 => "00000100000000011111101100000100",
9579 => "11111101000000000001000000000101",
9580 => "11111101111110111111111100000011",
9581 => "11111110000000110000000011111110",
9582 => "11111111000000000000001011111111",
9583 => "00000110111111110000010100000001",
9584 => "00000101000000100000001111111110",
9585 => "00000100111111110000011111111100",
9586 => "00000110000000011111111011111111",
9587 => "11111100111111110001100100000011",
9588 => "11111101000000110000001011111111",
9589 => "00000001000000001111111100000010",
9590 => "11111110000001010000001000000010",
9591 => "11110000111111100000010011111100",
9592 => "00001000111111001111111011111111",
9593 => "00000010000000010000010111111010",
9594 => "00000100000000111111110111111110",
9595 => "11111111111111110001011000000110",
9596 => "11111110111111011111110100000001",
9597 => "11101110111110011111100111110010",
9598 => "11110111111011011111111111111100",
9599 => "11111011111110101111110100000101",
9600 => "00000001111111001111001111111111",
9601 => "11101010000000111111111100001001",
9602 => "11111010111001111111100011111000",
9603 => "11111101111101111110110100000110",
9604 => "11110100111111101111100111110110",
9605 => "11110110111111000000100011111100",
9606 => "11101110111010001111110111110011",
9607 => "11110101111110101111101011111111",
9608 => "00001001111111001111000011111111",
9609 => "11111011111010000000011000000001",
9610 => "00000011110111101111110111101011",
9611 => "11110001111101111111101100000011",
9612 => "11110100111110011111000011101010",
9613 => "11101110111110100000010111111100",
9614 => "11100101110110011111100111110010",
9615 => "11110000111011111110011111110001",
9616 => "00000110111001011111000011111100",
9617 => "11110000110110000000111000001011",
9618 => "00001101110101100000100011011110",
9619 => "11110001111110110000001000000100",
9620 => "11101101111101101111001111101010",
9621 => "11101011000010000000001111110000",
9622 => "11011100110101011111001111101110",
9623 => "11100010110110111101101111100011",
9624 => "00001000110110101111000100000010",
9625 => "11101000111001001111110111111001",
9626 => "11111011111011111101010111101100",
9627 => "11111101111011001111110100000110",
9628 => "11100011111100011111100111011000",
9629 => "11110000111000000000011011110101",
9630 => "11001111111010111111101011110110",
9631 => "11111011111010111101011111111010",
9632 => "00000001110111111111001011111010",
9633 => "11101111111010011111110011111100",
9634 => "11111010111010100000001011001011",
9635 => "11110010111110111111011100001011",
9636 => "11110011111111011111011111011001",
9637 => "11101001111000110000010011111110",
9638 => "11001111110011101111111111110001",
9639 => "11011101111011011110011111101100",
9640 => "00000111111000101111011100000010",
9641 => "11101111110101011111100000000101",
9642 => "11111010110111001110100011010111",
9643 => "11111010111100101111101100000111",
9644 => "11110000111101001111111111100000",
9645 => "11110011111100001111100111111101",
9646 => "11011010101001110000010011110001",
9647 => "11100111111010011110100011100110",
9648 => "00000001111001011111000100000101",
9649 => "11111001110111100000010000000001",
9650 => "11111110110100111101101011011100",
9651 => "11110011111111010000000000000110",
9652 => "11101100111101101111001111100110",
9653 => "11100011111011000000101011110110",
9654 => "11011111101110001111110111111000",
9655 => "11010001110100111110101111100001",
9656 => "00000011101111001111001100000100",
9657 => "11110010110101111111101011110101",
9658 => "11110001110110101110100111100110",
9659 => "11110101111101011111111100001000",
9660 => "11101000111111011111001011100110",
9661 => "00000000111001011110100111110100",
9662 => "11101000000000011111101011110010",
9663 => "11101100111000011111101111110000",
9664 => "00000001111101001111010000001000",
9665 => "11011000111010111110110111101100",
9666 => "11100000111110101110000100010001",
9667 => "11110011111100011110101000000011",
9668 => "11111010111100111111000111111100",
9669 => "11110100111010111110100011101010",
9670 => "11101101000000011111101111110110",
9671 => "11000100111110111111100100000000",
9672 => "00000011111100001111010111111111",
9673 => "11111110111011011110100111110110",
9674 => "11011010111011001111110011111110",
9675 => "11110110111010101101110100000110",
9676 => "11110010111010011111010011111101",
9677 => "11110111110111111111001011010111",
9678 => "11110001111110011111110111110010",
9679 => "11011011111001110000010011110111",
9680 => "00000011111100011111100111111111",
9681 => "11100011111100001110011111101000",
9682 => "11010011111011011110100011111111",
9683 => "11011001111001101101001000001000",
9684 => "11110100111010001101111111111100",
9685 => "11110111110101111111011111110011",
9686 => "11110100000000111111101111110110",
9687 => "00000100111011100000000000000000",
9688 => "00000111111100111111101100000000",
9689 => "11110111110100001111110000000010",
9690 => "11011011000000001111100111111110",
9691 => "11101111111110001110010000001001",
9692 => "11111011111110001111011000000011",
9693 => "00010100000100010000101100010011",
9694 => "11110001000010111111111100001010",
9695 => "00001001000010011111110000000101",
9696 => "00000010000010100000110011111100",
9697 => "00010010000010010000101100001010",
9698 => "00010100000010010001011011111001",
9699 => "00000011000011110001100100001001",
9700 => "00010000000100000000000111110000",
9701 => "11111110000101100000001011111110",
9702 => "00010101000100011111010111111101",
9703 => "00000100111110000001001100000110",
9704 => "00001001111110111111101000010101",
9705 => "11101101000011111111110011111100",
9706 => "00000011000100001111101000010010",
9707 => "00001011111110101111100000000111",
9708 => "11111010111111001111010000010010",
9709 => "00001100000010100000100011111110",
9710 => "00001111000110001111101000000001",
9711 => "00000010000010110001000100000100",
9712 => "00001110000011110000000000001111",
9713 => "00000000111100000000101000000100",
9714 => "00011001000001100001000100010010",
9715 => "11111010000000111111110000000110",
9716 => "00001000000000001111111000010001",
9717 => "11110010000101011111010000000001",
9718 => "00010100000110100000001111111011",
9719 => "00000111000000010001100011111101",
9720 => "00010100000101100000011000010111",
9721 => "11110101111010100000100100000001",
9722 => "00001011000000110000010100011010",
9723 => "11110110111110010000000000000110",
9724 => "00000101111101101111101100010110",
9725 => "11111100000101111111100000000110",
9726 => "11111101000100011111011011110111",
9727 => "00000011000000000000001000001011",
9728 => "00001100111110111111110000010000",
9729 => "00001010111001110001010111111001",
9730 => "00011010000001000000011000010001",
9731 => "11111101111111010000010100001010",
9732 => "00000011111101101111101100000010",
9733 => "11111111111010111111011100000100",
9734 => "00010100000110000000101111111110",
9735 => "00000001000001000000111000000101",
9736 => "00000101111111111111110000010010",
9737 => "00000001110111010000110100000000",
9738 => "00001010000000010000000000010110",
9739 => "00000010111101010000011000000011",
9740 => "00001000111101111111001100001110",
9741 => "11111101111101101111011000000100",
9742 => "00011001111101100001111111111100",
9743 => "11100100111110110001100011100101",
9744 => "11111111111110101111101100010100",
9745 => "11110111110110000000111111111100",
9746 => "00001011111001111111100100010011",
9747 => "00000001111110100000010100010010",
9748 => "11111110111110101111001100010111",
9749 => "11111110111100101111011100000010",
9750 => "00001000111111000001000111111001",
9751 => "11100100111010110001001111101001",
9752 => "11111000000000010000000000001001",
9753 => "11111010111011010000001011111101",
9754 => "00000010111100111111010100000100",
9755 => "00000001000000100000000100001111",
9756 => "11111001111101101111111000001100",
9757 => "11111110111101011111010100001001",
9758 => "11111111111010010000000011111000",
9759 => "11100111111101000000001111101111",
9760 => "11111111111011011111001111111011",
9761 => "11111000111111010000101100000101",
9762 => "11111111111101011110110000000011",
9763 => "00000110000001010000011000001011",
9764 => "11110100111111111111001111111110",
9765 => "11100111111100111111100100000101",
9766 => "11100011111011110000000011111011",
9767 => "11110000111101101110001111110100",
9768 => "00000100111010101111011100001101",
9769 => "11101010000001110000101011111011",
9770 => "11111110111111001110110011110001",
9771 => "11110110111110100000100000001110",
9772 => "11110110000000111111101111100101",
9773 => "11100111111111110000001000000000",
9774 => "11000111110101111101100111111111",
9775 => "11110101111111111100010011111110",
9776 => "00000001110101101111001100001000",
9777 => "11111010111111110000000000001000",
9778 => "11111110111011001111101011100001",
9779 => "00000101111110001111101100000101",
9780 => "11111110111111001111101111101000",
9781 => "11101011111110011111010111101100",
9782 => "11001100111000001110111011110110",
9783 => "11100101111010101100010111111000",
9784 => "00001011111000001110111000000110",
9785 => "11100111111101101111111011111100",
9786 => "11111000111011001101110111110000",
9787 => "11101111111011001111101000001011",
9788 => "11101010111101101111010111100000",
9789 => "11110011110101111111011011101011",
9790 => "11010011111101101111101011110010",
9791 => "11111100111000111110000000000011",
9792 => "00000101111000101111011100000001",
9793 => "11110011110011011110100011111001",
9794 => "11010101111111011111001011111100",
9795 => "11100101111100101101111100000100",
9796 => "11110111111110001111001011100000",
9797 => "00000111000111100000100000000110",
9798 => "00000101000100010000101100010000",
9799 => "00000010000100100000110100000111",
9800 => "00000011000101000000011100000010",
9801 => "00000111000101100001011111111111",
9802 => "00011111000001000000110000001100",
9803 => "00001001000010100001101000000101",
9804 => "00001100000010000000100100000110",
9805 => "00001001000111011111101100010001",
9806 => "00000101000001011111101011111000",
9807 => "00000100000001100001001000000101",
9808 => "00001010111111100000010100001010",
9809 => "11110100000001110001001100001001",
9810 => "00101000000010000000010100001011",
9811 => "00000011000011000001000000000101",
9812 => "00000100000011111111011100000111",
9813 => "00001000111101110000010100001010",
9814 => "11111101000100111110111000001000",
9815 => "00000000000000000000101000000100",
9816 => "00010101000010100000011000011000",
9817 => "11111111110100000001101111111100",
9818 => "00100000111111110000011100001111",
9819 => "11101101000010110000110000001010",
9820 => "00001010000010100000101000010000",
9821 => "00000010000100000000011011111101",
9822 => "00000101000111001111011111111001",
9823 => "11110100000000000000111011111110",
9824 => "00101011000001100000110100011000",
9825 => "11111011110111010001100111100110",
9826 => "00101111000000010000100100010100",
9827 => "11110110000001110000111000000011",
9828 => "00001000111110001111111100011000",
9829 => "00001010000010010000100111111011",
9830 => "11111101000101111111000011111100",
9831 => "00000010000011000000110100000010",
9832 => "00111100000100100000100000110000",
9833 => "00001001110011010001010111110001",
9834 => "00101011000010010000100100010001",
9835 => "11111111000000010000001111111110",
9836 => "00000110111111010000000100010010",
9837 => "11111000111011110000011100000001",
9838 => "00000110000001111111100100000101",
9839 => "11111010000010010000101011101111",
9840 => "00100101000001000000100000010011",
9841 => "00001101110101010001010111101110",
9842 => "00100010111111101111111000001000",
9843 => "11111100111111100000010100000100",
9844 => "00001001000000100000001100001000",
9845 => "00001000110110110000101100001010",
9846 => "11111110111111010000010011111110",
9847 => "11100100000001000000001111101000",
9848 => "11110001111111100000101100001100",
9849 => "00000001111000110000111111101011",
9850 => "00010001111100011111000000000001",
9851 => "11111010000010100000010100011001",
9852 => "00000011111110111111111000001110",
9853 => "11111111111001000000000100010111",
9854 => "11111101111110101111111100000011",
9855 => "11101110000000110000000011110010",
9856 => "11100111111111010000010011111100",
9857 => "11110101111101000000010111111111",
9858 => "11111110111111111111010011111010",
9859 => "00000101111111110000011000011000",
9860 => "00000111111111101111110100000100",
9861 => "00000010111101110000011100010110",
9862 => "11111101111111010000001000001001",
9863 => "11101110000011001111010011110001",
9864 => "11100011000001100000011000000110",
9865 => "00000001000001010000010000001011",
9866 => "00000001000000001111101011111111",
9867 => "00001010000000000000101000000101",
9868 => "00001100000011110000111100000000",
9869 => "11111101000000010000001100000101",
9870 => "11100110111011001111001000000000",
9871 => "11111110000001011101111011101101",
9872 => "00000011111110111111111111110000",
9873 => "00000011000011110000010100000110",
9874 => "00000010111110111111011011100110",
9875 => "00000010111100110000001100001110",
9876 => "00000010111101111111011111101000",
9877 => "11110100111111010000001000000110",
9878 => "11101101110111111111101100000110",
9879 => "00011001111111101101110000001111",
9880 => "11110011111011001111110111101110",
9881 => "00000110000010001111100000100000",
9882 => "11111100000001001111010011010110",
9883 => "00000110000000111111101000000011",
9884 => "00000001000001111111111011100100",
9885 => "11101101000001011111001000001001",
9886 => "11110010110110001111111011111100",
9887 => "11110011111101111101101100000011",
9888 => "00001001111010101110101111111010",
9889 => "11111100000001110000001100010111",
9890 => "00000100111100001101011011010010",
9891 => "00000111111000010000000100001000",
9892 => "11111011111011001111110111100000",
9893 => "11101100111010001110111011111100",
9894 => "11010111111011111110101111110011",
9895 => "00001001111011111101100000001110",
9896 => "00000110110111011111001100000110",
9897 => "11110010111010010000010100000001",
9898 => "11110101111101111110111011011010",
9899 => "11101010111011011111111000000100",
9900 => "11110001111111101111010011011001",
9901 => "00000010000101000000100000000101",
9902 => "00001101111101100000110000000100",
9903 => "11110011000001100000110111111011",
9904 => "00000100000000000000100100001000",
9905 => "00001001000100110000010011111100",
9906 => "00011001111110010000100000000100",
9907 => "00000111000001010001101000000011",
9908 => "00001000000000110000101100001111",
9909 => "00010001111001010000110100000111",
9910 => "00000011000100010000100000000000",
9911 => "11111101000001110000100100001010",
9912 => "00000011000100110000110100001010",
9913 => "11111111111001010000010000000001",
9914 => "11111100000001000000001100010000",
9915 => "11110000000011110000111000000011",
9916 => "00001010000100001111110100001000",
9917 => "00001101111000110000110011110010",
9918 => "11110111000010111110110000000011",
9919 => "11110111000000000000001011110011",
9920 => "00011100000001010000110100001001",
9921 => "00000001110000100000100111100011",
9922 => "00011011111110011111100100000111",
9923 => "00000001111110100000000000001000",
9924 => "00001000111101110000010000000000",
9925 => "00000100111010000000101111110010",
9926 => "00001000000010001111111011111111",
9927 => "11110000000001110000110011101110",
9928 => "00100011111111010000000100011011",
9929 => "11111100111000010001100011101110",
9930 => "00110000111110011111101100001110",
9931 => "11111111000000011111011000000101",
9932 => "00001000111110111111111000010000",
9933 => "11111100110110101111111111111001",
9934 => "00000100000100010000000100000001",
9935 => "11100101111110000000111111100111",
9936 => "00101111000000100000001100011001",
9937 => "11111111110111010001101011100100",
9938 => "00011101111101101111110100001111",
9939 => "11111010111111011111110000001011",
9940 => "00000001111110011111111100001100",
9941 => "00000011111000001111111011111100",
9942 => "00000000000000010000001011111001",
9943 => "11101010000000000000100011011110",
9944 => "00001101000000110000010100001110",
9945 => "11111100111010100000011011001100",
9946 => "00001001111110101111001000000001",
9947 => "11111011111100001111010000101001",
9948 => "00001111111101011111101100001011",
9949 => "00000011110110100000000100000100",
9950 => "00000011000000000000010000000000",
9951 => "11110100111101010000100011101000",
9952 => "00001111111111010000111000000001",
9953 => "00000000111100010000011011011101",
9954 => "11111111111101101111011000001000",
9955 => "11110100111101011111001100110001",
9956 => "00001001111101000000001100001001",
9957 => "00010001111010010000011100001110",
9958 => "00001001000001011111110100001000",
9959 => "00001101111110000000011000000110",
9960 => "11010111000001000000111011111101",
9961 => "00000100111110111111101011111011",
9962 => "11111010000001100000000000001000",
9963 => "00001001000010101110110000100101",
9964 => "00000011000001100000100100001000",
9965 => "00010000000000100000010000010111",
9966 => "00000010000011001111111100001111",
9967 => "00001000000001000000000100000011",
9968 => "11011011000011110000111111110110",
9969 => "00001001000100000000100000000010",
9970 => "00000010000001010000111100010100",
9971 => "00001011000011100000001000000111",
9972 => "00001000000011110000100100000001",
9973 => "00000100000000110000000100010110",
9974 => "11111101111100110000010000000111",
9975 => "00001100000000101110001100000111",
9976 => "11110111111101100000010111100001",
9977 => "00000111000001100000100100011000",
9978 => "11110110000010011111010111101111",
9979 => "00000100000000100000001111111111",
9980 => "00000111000010000000001011101010",
9981 => "11111011000010101111111000001111",
9982 => "11110101111101011111101000000011",
9983 => "00000110000001001110000000001101",
9984 => "11111100111111110000010011011100",
9985 => "00000110000011001111111000001010",
9986 => "11110101000000101110101011100101",
9987 => "11111111111111110000100000000110",
9988 => "00001001111111110000001011100011",
9989 => "00000010000001001111111100000000",
9990 => "11111111111101010000011111111100",
9991 => "11100111000000001111101111110100",
9992 => "00000101111011100000001011100110",
9993 => "11110100000011111111111000001101",
9994 => "00000000111100111111011111101111",
9995 => "00000000000001000000010000000011",
9996 => "00000100111110011111110011101011",
9997 => "11110001111001001111011000000000",
9998 => "00000100111011110000011011111001",
9999 => "11111001111111011111011000001100",
10000 => "11111110111110101111011100000001",
10001 => "11101011111010101111001100000101",
10002 => "11011110111100111110000111111000",
10003 => "11100010111011001110100000000101",
10004 => "11110111111111111111111011111010",
10005 => "00010011000000110000101000001010",
10006 => "11110111000101010000000000000011",
10007 => "11111111000011001111110111111111",
10008 => "00000011000100010000011111110111",
10009 => "00001000000000010001011100001010",
10010 => "00010110111111000001001011111000",
10011 => "11111110000010100001111100000111",
10012 => "00010000000000000000010111111111",
10013 => "00000110110111110000100000001010",
10014 => "00001110000000000000011000001111",
10015 => "00000001000001010000110100000101",
10016 => "00001001000001100000110100000110",
10017 => "11111111111000000000111111111101",
10018 => "00001011000011001111111100001010",
10019 => "11110101000001100000111000000011",
10020 => "00000110000100010000010000010011",
10021 => "00000101111001110000110011111001",
10022 => "00000110000011000000100000000010",
10023 => "11101100000000110000001011101111",
10024 => "00000101000001000000100011111110",
10025 => "00001111111010101111111011101001",
10026 => "00000110111111111111101000000001",
10027 => "00000101000000011111110000000010",
10028 => "00000110000000110000001100001000",
10029 => "11110101110101011111110000000000",
10030 => "00001011111100010000111111111001",
10031 => "11110011000001101111111111110010",
10032 => "00001010000001101111111100001001",
10033 => "00000011111011000001110000000101",
10034 => "00001001111111001110101000000000",
10035 => "11111011111100001111100100001010",
10036 => "00000110111111001111110100001110",
10037 => "11110010111000001111001100000001",
10038 => "00010011111001010001100111110110",
10039 => "11101010000001000000101111100110",
10040 => "11111001111110000000001000000101",
10041 => "11110110000000010000011111101000",
10042 => "11111010111101001110001100000101",
10043 => "11111000111001101111000000010111",
10044 => "11111100111101111111100000010111",
10045 => "11110111111111101110110111110010",
10046 => "00000111111001100000111011110110",
10047 => "11100100111011100000011111011010",
10048 => "00010001111111000000100111111011",
10049 => "11111010000000111111010011010101",
10050 => "11101110111010111101100100000100",
10051 => "11110010110110101101101000101100",
10052 => "11111111111001101111011000000110",
10053 => "11111011000001101111110011110111",
10054 => "11111100111111111111111111111110",
10055 => "00010101111011010000000000010001",
10056 => "00000101111111100000011000000100",
10057 => "00000011000001101101001111011100",
10058 => "11010110000001111111110000001101",
10059 => "11111111111100111100001100100011",
10060 => "11111001111111010000001011111100",
10061 => "00000011000101100000010100001000",
10062 => "00000001000000000000111111111100",
10063 => "00011101111111111111110100011101",
10064 => "11100100000000010000000011111100",
10065 => "00001001000110101100111011111101",
10066 => "11110011000011011111101111111110",
10067 => "00001111111111001101100000000000",
10068 => "00000001000010110000011011111001",
10069 => "00001100000001100000101100001000",
10070 => "00001000000010000000101000010001",
10071 => "00010001000010011111101000001100",
10072 => "11010011000001010000110011101010",
10073 => "00001001000100001110011111111001",
10074 => "11110110000100000000000000000101",
10075 => "00000111000001111111111100000100",
10076 => "00001001000010000000010111110101",
10077 => "00001001000000110000001100000100",
10078 => "00001010000001010001000011111010",
10079 => "11101100000010101111010011101101",
10080 => "11110011000010010000010111101010",
10081 => "00000000000100101111110111111011",
10082 => "11101111111110101111100111111011",
10083 => "00000000000000001111110100000000",
10084 => "00000111000000101111111100000010",
10085 => "00000111000010110000000100000110",
10086 => "00000010000001000001000000000110",
10087 => "11111011000000011111001000000010",
10088 => "11111100111111100000011111111011",
10089 => "11111011000100101111111100001110",
10090 => "11111110000001111111010111111111",
10091 => "00000010111111101111100100000010",
10092 => "00000110111111100000100011111000",
10093 => "00000101000000100000000111110101",
10094 => "00000100111101110000000111110101",
10095 => "11011011000000011110110111100000",
10096 => "11111111000000111111111011101111",
10097 => "11110000000000100000011100001000",
10098 => "00000001111000101111011011100101",
10099 => "11101111111111001111101100000011",
10100 => "11111010111110001111000011110101",
10101 => "11111010111010011111110100000011",
10102 => "11111111111011101111101111110100",
10103 => "11101101111101111111011011111000",
10104 => "00000110111110011111100100001000",
10105 => "11101111111001110001000000010110",
10106 => "11110111111101001111001000000010",
10107 => "11111011000000000000011000000111",
10108 => "11110101111110101111001011111111",
10109 => "00010000000001000000111000010000",
10110 => "00010100000100110000010000001110",
10111 => "00001010000100000001001100001001",
10112 => "00000011000010110001000000001110",
10113 => "00010000000001000000101000001100",
10114 => "11111110000011110001100000001100",
10115 => "00000101000010110001110000000110",
10116 => "00001011000011100000111000010000",
10117 => "11111010111010110000010100000001",
10118 => "00011110111101000001111100001100",
10119 => "00001001111111110001000100000111",
10120 => "00000100111111100000010000001100",
10121 => "00001000000001001111111100000110",
10122 => "11101111000010111111000000001010",
10123 => "00000100111110011111011100000011",
10124 => "11111110000010000000101000010011",
10125 => "11111000111000110000110000000000",
10126 => "11111111111011000000111100000011",
10127 => "11111111000011101111011111110111",
10128 => "11111010000001100000010011110101",
10129 => "00001010111111001111111011111011",
10130 => "11101010000000011111110111110111",
10131 => "00000000111100011111001000000100",
10132 => "00000110111111110000001011111100",
10133 => "11111010111000001111110011110100",
10134 => "00010000111000010001110111111010",
10135 => "11110100111101000000111011101011",
10136 => "00001101111110000000000000001011",
10137 => "11111100000001110000010000010000",
10138 => "11100000111110101110110111111110",
10139 => "11111010111100011110010000010110",
10140 => "11111010111101001111001000001101",
10141 => "11101110111100101111010100000010",
10142 => "00010111110110100011000011101111",
10143 => "00001011111101110001110000001010",
10144 => "00001010111100011111011000000111",
10145 => "11110101000101110001001000110010",
10146 => "11101101111100101110110000000011",
10147 => "11110100111011011111001100101100",
10148 => "11110111111011101110110000010000",
10149 => "11110010000000111110101011111110",
10150 => "00000011110101100010010111110000",
10151 => "11110110111001101111111111111100",
10152 => "00001011111011001110111011011111",
10153 => "11101001000111110000011000010101",
10154 => "11101010111010001101011111110001",
10155 => "11100111111000101110111000110101",
10156 => "11110011111011011111010011110010",
10157 => "11100100111101011111100011110101",
10158 => "11011001111010101111100011111000",
10159 => "00011010111010011101110000011101",
10160 => "00000011111010001111010011111001",
10161 => "11110110111110111101001011101100",
10162 => "10111100000001101110100011101000",
10163 => "11100111111010001101111100010011",
10164 => "11110010111100101111101011101000",
10165 => "11110110111101110000000011111111",
10166 => "00000001111011110001001100000100",
10167 => "00011001111100101111101000011000",
10168 => "11111100111101000000010100001101",
10169 => "11111110000000101011010100000001",
10170 => "11101010000011101111101111110111",
10171 => "11111111000000101111001100011111",
10172 => "11111111111111110000001000000000",
10173 => "00000110111111100000011100000001",
10174 => "00001011000000110000011000000100",
10175 => "00000110111111100000001100000000",
10176 => "11110111000010010000001011110011",
10177 => "00000111111111001111101100001101",
10178 => "00000001000000100000010111111111",
10179 => "00001000000010111111111100001001",
10180 => "11111111000010000000000100000100",
10181 => "00010000000010010001010011111001",
10182 => "00000111000010010001000100000001",
10183 => "11111111000001001111110111111111",
10184 => "00001000000011110000011111111100",
10185 => "00001011000011110000111100000111",
10186 => "00010011111111000000111011111111",
10187 => "11111011000100100000000100001101",
10188 => "00000010000010100000100000000100",
10189 => "00000010000010000000110100000000",
10190 => "11110011000010011111101000000001",
10191 => "11111001000100011110111000000100",
10192 => "00000001000001010000001100010110",
10193 => "00001000000001000000100100001100",
10194 => "00010010111111110000011011111010",
10195 => "00001010000011100000001011111100",
10196 => "00000011111111111111110111111110",
10197 => "11110000000000110000101011111011",
10198 => "11101111111010011111100011110110",
10199 => "11100111000001001110111011101110",
10200 => "00010010111001011111100000011001",
10201 => "00000010000000000000100000000001",
10202 => "00001001111101101111011111111111",
10203 => "00001101111011000000010100000110",
10204 => "11111000111101111111111111110001",
10205 => "00000100111101000000001111100000",
10206 => "00001101111110010000110111110101",
10207 => "11110101000011000000110111111110",
10208 => "11111111000101011111101100010100",
10209 => "11111010111101001111001111100011",
10210 => "11110110000000100001110000010101",
10211 => "11100000000011101110100000000110",
10212 => "11110110111101001111000100010001",
10213 => "00001001000001000000001100000101",
10214 => "00010100000011010000010100000010",
10215 => "00000000000001000001100000000001",
10216 => "00001010000000010000000100001101",
10217 => "00001000000001010000000100000110",
10218 => "11111111000001000000010000010001",
10219 => "00000011000000100001011000001000",
10220 => "00000100000001010000011100011011",
10221 => "11110010111101111111101100000111",
10222 => "11111111111100000001010000000010",
10223 => "00000111000000001111111100000100",
10224 => "11111101111111010000000100000001",
10225 => "00000010000101111111110100000010",
10226 => "11011100000001001110111011111110",
10227 => "00000101111110110000110000001010",
10228 => "11111000000000110000011111111011",
10229 => "11101111111010010000000011111010",
10230 => "11111000110111000001101000000010",
10231 => "00000101111111001111101100000110",
10232 => "11110001111010110000000011101100",
10233 => "00000011001000101111011100010000",
10234 => "11001110000000011111010111101010",
10235 => "11111111111100001110100000001011",
10236 => "11111001111111001111110111110001",
10237 => "11101011111101111110011100000010",
10238 => "00000111111000010010010011110110",
10239 => "00010011111110101111110100001100",
10240 => "11110110111011011111100111110000",
10241 => "11111011001101111111110000110001",
10242 => "11001010000001001110111111101100",
10243 => "11111010111100101110110000001100",
10244 => "11110111111101101111000111111000",
10245 => "11101100000001111110100000001001",
10246 => "00011000110110010011110011110100",
10247 => "00010110111100000000100100011110",
10248 => "00000001111011011111011011110011",
10249 => "11101100001111110000110100111111",
10250 => "11101010111110011110011011110101",
10251 => "11110111111010110000011100100011",
10252 => "11110100111010111110110100000110",
10253 => "11110011111100011111000011110011",
10254 => "11110011111000110000100111101110",
10255 => "11111110111010111110011100001000",
10256 => "00000001111011101111001111011011",
10257 => "11101011000101111111010111110110",
10258 => "11011101111101001110010111101011",
10259 => "11101100111001111111000100101100",
10260 => "11110011111100001111010111101001",
10261 => "11110011110111101111111011111100",
10262 => "11011100111110111100100111110101",
10263 => "00001100111100111100000100001011",
10264 => "00010110111101011111110111100111",
10265 => "11101110110010111101101011100111",
10266 => "11000111000001111110110111011001",
10267 => "11101010111111011110101000110110",
10268 => "11111010111111101111000111100011",
10269 => "00000000111100110000101100000011",
10270 => "11111101000000101111111111111110",
10271 => "00010010000010001111100100010111",
10272 => "00010111111111010000001011110000",
10273 => "00000001111101011110101111110100",
10274 => "11110101000001110000010011110011",
10275 => "11110111000000111111101000100110",
10276 => "00000010000001010000000011111001",
10277 => "00000011111110100000100000000111",
10278 => "00001100111111110000111100001000",
10279 => "00000111000011110000101000010000",
10280 => "00000111000001010000010000001000",
10281 => "00000100111111011111111100000001",
10282 => "00000001000011001111011100000111",
10283 => "00000111000001110000100100000001",
10284 => "00000011111110110000011100010110",
10285 => "00001011000011010000101100000011",
10286 => "00001011000011100001010100001101",
10287 => "00010111000011010000101100010010",
10288 => "00001010000001000000001000000100",
10289 => "00000010000010000000001000001110",
10290 => "00000011000011111111110000001001",
10291 => "00000011000001010000001000001011",
10292 => "00001010111111110000011100001101",
10293 => "11111000000010010000101000000001",
10294 => "00000000111101110000001011111110",
10295 => "00000110111110101111010000000010",
10296 => "11111111111110000000000111111101",
10297 => "00000000000011001111101011111110",
10298 => "00000001111111111110011011110011",
10299 => "00010001111110011111100100000100",
10300 => "00000100111111000000011111111010",
10301 => "11111000000010110000001000000100",
10302 => "11110011111001110000010111110100",
10303 => "11101011111100001111001011111111",
10304 => "11111010111110001111011011110100",
10305 => "00000011000100001110111000000101",
10306 => "00000000111011101111001111110000",
10307 => "00010000111010101110110100000101",
10308 => "11110011111110011111100111111000",
10309 => "11100011111011101110011011100110",
10310 => "11010110110101011110101011101010",
10311 => "11101110110100011101111011111011",
10312 => "00001000110101001110010100000000",
10313 => "11101001111001110000000100001010",
10314 => "11101111111011011101101111100011",
10315 => "11010010110111101110111000001001",
10316 => "11100000111011011110100111011110",
10317 => "11111111000100101111100111111011",
10318 => "11111000111110111111101111111100",
10319 => "11101011111111000000001011110101",
10320 => "00000110111110011111100111111100",
10321 => "00000001000011110000100100000101",
10322 => "00010110111011001111110011110001",
10323 => "00000011111111110001010000000100",
10324 => "11111011111110101111110111101010",
10325 => "11111101000001100000101111111011",
10326 => "00000000111100000000000000001000",
10327 => "11111100111111011111010011111101",
10328 => "11111010111100100000001100000000",
10329 => "00010101000100111111111111101101",
10330 => "00000001111111100000011111111011",
10331 => "00000100111110011111010100000011",
10332 => "11111001000000010000011111111100",
10333 => "11111000000001011111001011111010",
10334 => "00000001110111100000110111110000",
10335 => "11111001111100111111110111111100",
10336 => "00000010111011001111111011111001",
10337 => "00000001001000011111110100001100",
10338 => "11101010111110101110111011101001",
10339 => "11111110111011011110101000001110",
10340 => "11110100111100111111001111110001",
10341 => "00000000000111111111101011111010",
10342 => "00000110111000010001110011111001",
10343 => "00010010111100110000011000001111",
10344 => "00000110111110001111010100000011",
10345 => "11111111001100111111100000101111",
10346 => "11101110000000011111100100000011",
10347 => "11111100000000001111100000010100",
10348 => "11101101111111001110111100000011",
10349 => "11110010000110101111000100000011",
10350 => "00000000110100110001011011110110",
10351 => "00001000111011111111101100010000",
10352 => "00001000111100011111010111111001",
10353 => "11101100010000101111101000100110",
10354 => "11101011111110001110000011110010",
10355 => "11111111111101010000001100011111",
10356 => "11101010111110011111011011111110",
10357 => "11101111111111001111000100000011",
10358 => "11110110111101111110101111110101",
10359 => "00000010111101111110010000001100",
10360 => "00011011111101111111010111101001",
10361 => "11110001111110111111010111111111",
10362 => "11011101111110111110011111101111",
10363 => "11111110111110101111110000100101",
10364 => "11110101111111101111011011110100",
10365 => "11111100111110011111101000000010",
10366 => "11110101111111111110111100000111",
10367 => "00000011000000001111010000000100",
10368 => "00001110000000011111100011111110",
10369 => "11111001111011111110101011101010",
10370 => "11101011000010001111100111111101",
10371 => "11101011111101110000000000011111",
10372 => "11111001000000001111100000000110",
10373 => "00001011000001000000011111111101",
10374 => "00000000000001001111110100001011",
10375 => "11110111111111001110111111111111",
10376 => "00001000111111010000110111101011",
10377 => "00001011111111111100001011110100",
10378 => "11100101111110100000100111110110",
10379 => "11111100000010101110101100100110",
10380 => "00000110000000100000010111110111",
10381 => "11111110111111100000011000000011",
10382 => "00001101000010100001000111111101",
10383 => "11101110000001100000001011101111",
10384 => "00000011000010100000001011101000",
10385 => "00000101000000110000101100100111",
10386 => "11111000111011101111100011111011",
10387 => "00000100000001001111110100000110",
10388 => "00001010111101100000011100000010",
10389 => "00000010000001000000011100001110",
10390 => "00010110111111100001100100000101",
10391 => "00000011000100100000110011111110",
10392 => "00001110000001100000011011110110",
10393 => "11111101000010010001011000101011",
10394 => "00000000111111001110111000000011",
10395 => "11111001000000000001011100000100",
10396 => "00001011111110100000100000000110",
10397 => "11111100000010010000000100000011",
10398 => "00000111111101100001101000000100",
10399 => "11011010000000110000001011100011",
10400 => "11111100111111111111110111110001",
10401 => "11111001000011110000000000001101",
10402 => "00000011111011101110100100000001",
10403 => "00000100111100011111111000001001",
10404 => "00000111111100100000000000000011",
10405 => "11111101000000011111001111111011",
10406 => "00000101111101110000000011110110",
10407 => "00000010111110110000010100000101",
10408 => "00000010111101101111110100000000",
10409 => "11101100111111101111011011111001",
10410 => "11111000111100011111101100000010",
10411 => "11110110111010101111001000000011",
10412 => "00000011111101011111011000000101",
10413 => "11011011111110111101100011110010",
10414 => "11101100110110011111101011101111",
10415 => "11111010000000101111001100000010",
10416 => "00000110111100101110110011111110",
10417 => "11100111111100100001011011111101",
10418 => "00010000111100101100110011110100",
10419 => "11010010110100111111111000000011",
10420 => "11111101111011001111001011101110",
10421 => "11111011000101101111110111110111",
10422 => "11111010111110000000110111111001",
10423 => "11100100000010001111111111110000",
10424 => "00001000111111101111111011111100",
10425 => "00000100000100110000111000000010",
10426 => "00010001111010011111011011110101",
10427 => "00000000111110110000011000001001",
10428 => "11111011111101010000000111111000",
10429 => "00000000111101011111101100000100",
10430 => "11111101111111000001000011111110",
10431 => "11111100111101010000000011111101",
10432 => "00001100111110001111101000000000",
10433 => "00000000111110111111110011111111",
10434 => "11110010111111001111111011110111",
10435 => "00000100000000001111011000000011",
10436 => "11110011000001011111101111110101",
10437 => "11110010111111101111100011110100",
10438 => "11110001111001110000100111111101",
10439 => "11111001000000011111001111110110",
10440 => "11111101111001111111011011110000",
10441 => "11110100000011101110100111111111",
10442 => "11011000111101111111010011101011",
10443 => "11110110111100001110110000001010",
10444 => "11111001111100111111111111110001",
10445 => "11110100111110011110111011110000",
10446 => "11110010111100100000010011110111",
10447 => "11110100000000111111001011111010",
10448 => "00001011111101011111110111111000",
10449 => "11110000111111001110100100000000",
10450 => "11010100111011101110101011101100",
10451 => "11111001111010001110110100001011",
10452 => "11111100111100011111011011110011",
10453 => "11110111000001101111000111111001",
10454 => "11111001111100110000100011110101",
10455 => "11111000111110001111010111111100",
10456 => "00000101111101011110111111110010",
10457 => "11110100000010011111001000001111",
10458 => "11100000111110111111100111101000",
10459 => "11110010111110101111101000010010",
10460 => "11110010000001001111100011101111",
10461 => "11111011000011000000000000000001",
10462 => "11110000111100101111110111111010",
10463 => "00001100111110101110010000001111",
10464 => "11111011111110011111110111101010",
10465 => "11111001000010111110110011111111",
10466 => "11100110000000111111111111101001",
10467 => "00000011111111011111110000010010",
10468 => "11111000000010101111111111101010",
10469 => "00001000000100000000100000000100",
10470 => "11110110111111100000000000000001",
10471 => "00010000111111001110110000001010",
10472 => "00001110000000010000010011100110",
10473 => "00001000000011011110010111110100",
10474 => "11111001000001110000000011110110",
10475 => "11111101000000011110111100011011",
10476 => "11111011000001000000010011100111",
10477 => "00001100111111110000011011111001",
10478 => "11111001000001101111011000000000",
10479 => "00001010111101111111001000001001",
10480 => "11110100111111111111111100000100",
10481 => "00001000000000111011100111111110",
10482 => "11100111000001000000011111111110",
10483 => "00001100000000001101100100001010",
10484 => "11111001000010100000100011110111",
10485 => "11111110111111010000100011111100",
10486 => "11111111000000101111111111111111",
10487 => "11110100111110011111110011111110",
10488 => "00000101111100101111110000000011",
10489 => "00000010000000001101101011111101",
10490 => "11100010111011101111101111111111",
10491 => "11111110000000101110100000001111",
10492 => "11111110000000010000010011111110",
10493 => "11110100111111111111111011110110",
10494 => "00000010111100100001000011111000",
10495 => "11101101111111100000100111110100",
10496 => "00000001111101101111100111111010",
10497 => "11111000000000011111011111111100",
10498 => "11100100111101101111000000000010",
10499 => "11111110111011001110110100001101",
10500 => "00000000111010111111110011111101",
10501 => "11111101111111001111111011110011",
10502 => "11111011111100000001000011101011",
10503 => "11010001111100111111111111011110",
10504 => "00000001111100111111101011101110",
10505 => "11110110000000111111010100010100",
10506 => "11100010111000001110100011110100",
10507 => "11111001111011101110100000001100",
10508 => "11110111111010011111101011101111",
10509 => "11110000111010111111010111110010",
10510 => "11101110111010111111100011110010",
10511 => "00001011111001111111101000000111",
10512 => "00000101111000101111010100001101",
10513 => "11101010111011101111001000001110",
10514 => "11101011000000001110100011111010",
10515 => "11100100111101011110001100001000",
10516 => "11111000111101001111010111101110",
10517 => "11101000111110011110111111110001",
10518 => "11111111110111010000111111111011",
10519 => "11111110000001110000011000000000",
10520 => "00000111111100111111001100010011",
10521 => "11110011111101110000101000000001",
10522 => "00001000111101111110000000000010",
10523 => "11101010111010001111101100000100",
10524 => "11110111111101001111100011111100",
10525 => "11110000000000111111100011110000",
10526 => "11011001111110000000000011110100",
10527 => "11011100111101011101111011100011",
10528 => "00000010111100101111001111110110",
10529 => "11111011000000000000010011110011",
10530 => "00000000111000011111011111011110",
10531 => "11111010111100010000111000000111",
10532 => "11111000111100011111000111010011",
10533 => "11111000111110010000000100000001",
10534 => "11110110000000111111000111110110",
10535 => "11111101000000001111100100000001",
10536 => "00000011111111111111100100000010",
10537 => "00000100000000000000000100000011",
10538 => "11111001111111010000001111111000",
10539 => "11110010111110000000001000001000",
10540 => "11111000111111111111101111111100",
10541 => "00000010111101011111110100000111",
10542 => "11101100000000111111111111111101",
10543 => "11111110111111111111001000000101",
10544 => "00000111000001010000000111110000",
10545 => "11110111000000010000010000010101",
10546 => "11101100111110110000010111100101",
10547 => "11101110000100100000100000000101",
10548 => "11111110000001011111011111101111",
10549 => "11110000000011001110111100001010",
10550 => "11111101111100100000000000000010",
10551 => "11111110111101001110011011111010",
10552 => "00000111111010011110111111011111",
10553 => "11100111000000001111110000100000",
10554 => "10111111111111101110111111011011",
10555 => "11111100000000100000111000001100",
10556 => "11110110000001011111111111101010",
10557 => "11101110000110101111101100001000",
10558 => "11111001111010100000101000000000",
10559 => "00001100111111011110000100000110",
10560 => "11111011111101011111010011001110",
10561 => "11101001000110011110110000001111",
10562 => "10110011111111011110100111100001",
10563 => "00000011111110010000100000001101",
10564 => "11110011000001011111111111100111",
10565 => "00000001001001010000001111111110",
10566 => "11101101111110110000000011111110",
10567 => "00001001000000111101111000001101",
10568 => "11110110111101101111100011100110",
10569 => "11111110000110011101010011111110",
10570 => "11101001000001001111110011100011",
10571 => "00000100000000011111100000001001",
10572 => "11111011000001100000000011100110",
10573 => "00001000000101000000011011111011",
10574 => "11101100111100101111010100000101",
10575 => "00001000111111111110011100010001",
10576 => "11111100111110000000000011111011",
10577 => "00000011000011011100101011110111",
10578 => "00000011000000110000001111110111",
10579 => "00000001000001001111011000001010",
10580 => "11111000000001000000010011101110",
10581 => "11111001000010011111111011110011",
10582 => "11101001000000111101110100000000",
10583 => "00001011000000011101010000001111",
10584 => "00010001111101110000000100010100",
10585 => "00000010111111011101101011101110",
10586 => "00000001000000110000010011110001",
10587 => "11111111000001001101100000010100",
10588 => "11111111111111000000001011101111",
10589 => "11111111000000110000000011110011",
10590 => "11110000000001001110111011110000",
10591 => "00000110000000001110001000001010",
10592 => "00001000000000001111101100001010",
10593 => "00000001111111101110011111011110",
10594 => "11111110000000010000100011111000",
10595 => "00000111111111111101011100001011",
10596 => "11111101111111011111010111110011",
10597 => "11111001111111011111011011100110",
10598 => "11110100111101101111010011110001",
10599 => "11101001111101001111000011101011",
10600 => "00000111111100011111000100000001",
10601 => "11111100111110111110000011010000",
10602 => "11111001111100101111011111110000",
10603 => "11111001111011101101000100000011",
10604 => "11111111111011101111011111101111",
10605 => "11110000111111111111010111110000",
10606 => "11110010111010111111100111101110",
10607 => "11101100111111101111000111111011",
10608 => "11111110111101111110110111111111",
10609 => "11111101111101111110100000000000",
10610 => "11110111111011111111110011111011",
10611 => "11111100111100101101011100000101",
10612 => "11110111111100011111000011110110",
10613 => "11011111111010001110011111110100",
10614 => "11100110110111011110110011101101",
10615 => "11111110111100001110101111110100",
10616 => "00000101111000011110011100001000",
10617 => "11100001111010111110001011110101",
10618 => "11101001111110011101101011101011",
10619 => "11011101111000111101000000000110",
10620 => "11100100111010101110110111100110",
10621 => "11101101111110011110111100000000",
10622 => "11111010111100100000010111111001",
10623 => "00000001000000111111100111111110",
10624 => "00001001111100111111110111111110",
10625 => "11110110111110011111101100001101",
10626 => "11110010111111011110011111110101",
10627 => "11110101111001101111111100000011",
10628 => "11111010111101111111100111101010",
10629 => "11111010000001100000000011111100",
10630 => "11110000000001001111110111111001",
10631 => "11110111000001111110100011110101",
10632 => "00000110111111001111111011111001",
10633 => "11111011000000110000111000000100",
10634 => "00010100111100010000001111110010",
10635 => "00000010111111110001000000001001",
10636 => "00000000111101111111110111110011",
10637 => "00000000000000010000000100010111",
10638 => "11110111000110101111011100001000",
10639 => "11111101000011001111110000000010",
10640 => "11111110000001000000011011111100",
10641 => "00000011111010000000110100001111",
10642 => "00000111111111100000111111111100",
10643 => "11111100000101100010101000000000",
10644 => "00001001000011110000001011111001",
10645 => "11111111000010001111100000010011",
10646 => "00000000000010101111111100000100",
10647 => "00001011000010111111110000001111",
10648 => "11111000000001000000001111111010",
10649 => "00001000000011001110100000001100",
10650 => "11010101000010111111111011111011",
10651 => "00010010000001000000110000000010",
10652 => "00000011000011000000111111111011",
10653 => "11110100001011011110111011111110",
10654 => "11110110111101110000111000001001",
10655 => "00000000111111011110110100001000",
10656 => "11110001111111001111110111011101",
10657 => "11111111001000001101100100000001",
10658 => "10111010111111101111010011101100",
10659 => "00001110111111011111100100001101",
10660 => "00000011111110010000001011101101",
10661 => "11111000000110111111100000000011",
10662 => "11101111111100011111011111111100",
10663 => "00010010111110001110100000010101",
10664 => "11111010111101101111101111100100",
10665 => "11110111000100011100100011111010",
10666 => "10101101000010011110111011101011",
10667 => "11111110111111011110101100001000",
10668 => "11111110111111111111100011101100",
10669 => "00000110000110100000010111111010",
10670 => "11101011000001001110101000000101",
10671 => "00001010000001011110100000001001",
10672 => "00000111111101111111100000000001",
10673 => "11111111000011101010111111110011",
10674 => "11010010000010000000101011101110",
10675 => "00001011000000101110000000010011",
10676 => "11111011000000110000000111110011",
10677 => "00000001000101101111110111110011",
10678 => "11111000111011011111011000000100",
10679 => "00010110000000111111000000011100",
10680 => "00010110111111000000001100010101",
10681 => "00000001000100001101000111100110",
10682 => "00000011000100000000000011111111",
10683 => "00000000000001101101101100000100",
10684 => "11110101000011011111111011111010",
10685 => "00000100000110000000010111101010",
10686 => "11110001000000111111010011111110",
10687 => "00010111111110001111000000011000",
10688 => "00001101111101110000000100011000",
10689 => "00001100000010101100001111010000",
10690 => "11111101000011100001001111111010",
10691 => "00001011000000101011110000001100",
10692 => "11111011000000101111111111110110",
10693 => "11110110000011001111111111100110",
10694 => "11101110111111111111000100000001",
10695 => "00001100111100011110001100010011",
10696 => "00001000111011100000011000001100",
10697 => "00000110000010111100100011101001",
10698 => "11101110000001000000010111110010",
10699 => "00000010000000001100010100001111",
10700 => "11110111000000001111111011101001",
10701 => "11110101111111110000010011101001",
10702 => "11101011111111111110110111111011",
10703 => "11110100111000001101110111111110",
10704 => "00000111111010011111111011111111",
10705 => "00000111111101001110101111011011",
10706 => "00000001111101011111110011101000",
10707 => "11111111111111111110000000000111",
10708 => "11111100111101111111101111100100",
10709 => "11110010111111011111001111101100",
10710 => "11101001111101011111011011110001",
10711 => "11111110111110001110011000001000",
10712 => "00000101111110001111000011111010",
10713 => "00000010111110010000001111100011",
10714 => "00000001111101111111011111100111",
10715 => "00000001111010110000001000001011",
10716 => "11101101111111001110111011101100",
10717 => "11101001111011001110110111111000",
10718 => "11011111111001011110100111110100",
10719 => "00000011111010111101100100000001",
10720 => "00000010111001011111000011111010",
10721 => "11100010111010011110111111101110",
10722 => "11110001111110111101101111100101",
10723 => "11011010111010111110001000001011",
10724 => "11110010111101111110110011100001",
10725 => "11111010111100011111111000000011",
10726 => "11110100000000001111110011111100",
10727 => "00000111111110011111011100000101",
10728 => "00000100111111001111101100000000",
10729 => "11111111111001110000000111111111",
10730 => "11110010000000101111111011111100",
10731 => "11111110111111100000100000001000",
10732 => "11111001000000011111101011111011",
10733 => "00000001000001100000010100000010",
10734 => "00001000000000010000100000000010",
10735 => "00010000000000110000100100001001",
10736 => "00000001000001110000001100001010",
10737 => "00000110000000110000011000000011",
10738 => "00000100000100000000011000001110",
10739 => "00000011000000110010000000001010",
10740 => "00000010000000110000001100010110",
10741 => "00000100000010000001000011101101",
10742 => "00000011111101010001110000000010",
10743 => "11101101000001110000111011111011",
10744 => "00001010000001100000100000000001",
10745 => "00000100000011101111111011100110",
10746 => "00000000111101011111001000000101",
10747 => "00001100111011011111101100001001",
10748 => "11111001111101010000101000000100",
10749 => "00010011000001000001010111110000",
10750 => "00001010111101100000100011111110",
10751 => "11111111111111110001000011111000",
10752 => "00000111000001110000100100001011",
10753 => "00010000000010011110100100010001",
10754 => "11011010000010010001001100001000",
10755 => "00000111000100101110110000000110",
10756 => "11111000000010010000100100000111",
10757 => "00000100000110100000110000010100",
10758 => "00000100111110110000001100001010",
10759 => "00001110000000011111110100001110",
10760 => "11111000000001110000011111111111",
10761 => "00000101000111001110010000101101",
10762 => "11011101000001000001001000000000",
10763 => "00001011000110111111101100001101",
10764 => "11111111000110010000000100000011",
10765 => "11110110001001001111000100001010",
10766 => "11111110111110001111110000000100",
10767 => "00010000111110001111100000010010",
10768 => "00000100111111000000100111111000",
10769 => "00000011000011001110111000010101",
10770 => "11011001000001011111011011111010",
10771 => "00000110111110010001010100000011",
10772 => "11111001000010000000111011111111",
10773 => "00000010000100110000000000000000",
10774 => "11111011111111111111100000000101",
10775 => "00010000111100111111010100010101",
10776 => "00000110000000001111100100000100",
10777 => "00001011000011001110100111110110",
10778 => "11101101000001000000011111111000",
10779 => "00001100000001111111101100010000",
10780 => "11111110000100000000101111110101",
10781 => "11111100000011111111111000010001",
10782 => "11111100000001100000000100001010",
10783 => "00010110111101011111100100011010",
10784 => "00001010111110111111111111111110",
10785 => "00010010000001111111010000001011",
10786 => "00001100000010110000010011111100",
10787 => "00001001000001000000100000000011",
10788 => "00000011000001010000100111111011",
10789 => "00001000000110010000000100000011",
10790 => "11111000000010101111100000010000",
10791 => "00010101111110001111100000010011",
10792 => "00010100000000111111101000000111",
10793 => "00001011000001111111000000011010",
10794 => "11111110000011110000110000000010",
10795 => "00001100000010001111111100001011",
10796 => "11111111000001100000001011111101",
10797 => "11111111000001101111100000000011",
10798 => "11111000111110011111010000000000",
10799 => "00010011111110001111000100010110",
10800 => "00001011111111001111110111111111",
10801 => "00000101111110101111011000000110",
10802 => "11111010000011001111110011110100",
10803 => "11111101111111011110010000000111",
10804 => "00000000000010111111111111111111",
10805 => "11111111000001101111101000000101",
10806 => "11111101000001000000001111111111",
10807 => "11111111111110011111100100000001",
10808 => "00000111000001100000100011111101",
10809 => "11111101000000100001001000000011",
10810 => "00001000111101000000000111111010",
10811 => "11111111000000110000101000000100",
10812 => "00001001000000101111110111111100",
10813 => "11111111000001101111111011111111",
10814 => "11101011000001111111100100000000",
10815 => "00001000111110011110110000010100",
10816 => "00000110111101001111101111111100",
10817 => "00001011000000010000011100000010",
10818 => "00001100000000100000110011110100",
10819 => "00001100000010000000111000000001",
10820 => "00000010000000101111100111110001",
10821 => "11101100000010001111000100000000",
10822 => "11101000111011001110111111111100",
10823 => "00000110111110001101111000000001",
10824 => "00000101111111101111100011111011",
10825 => "11101110111111100001101011110010",
10826 => "00010110111111011110000111101101",
10827 => "11110001111110000010000100000110",
10828 => "11111100111101001111101111100001",
10829 => "11111110111110000000000111111111",
10830 => "11110011000000001111101100000010",
10831 => "00001000000000101111001000000011",
10832 => "00000100111111001111111100000001",
10833 => "00000001111011100000001011111011",
10834 => "11111010000000001111111100000001",
10835 => "11111011111110100001100000001000",
10836 => "11111111111111011111110011111001",
10837 => "00000000000000000000000000000000",
10838 => "00000000000000000000000000000000",
10839 => "00000000000000000000000000000000",
10840 => "00000000000000000000000111111010",
10841 => "11111101000000100000000000000011",
10842 => "11110011111110111111101111111101",
10843 => "11111001000000100000000011111110",
10844 => "00000001000000001111100100000011",
10845 => "11111010111111111111111111111000",
10846 => "11111101111110101111001011110110",
10847 => "11111010111111010000000111111101",
10848 => "00000010111110110000001011111101",
10849 => "11111110111110110000000111111101",
10850 => "11110110111111011111111011111001",
10851 => "11111001000000011111111111111110",
10852 => "11111011111111001111110000000000",
10853 => "11110111111111011111110111111100",
10854 => "11111011000000001111000011110101",
10855 => "11111111111110100000000111111110",
10856 => "11111010000000001111011111110010",
10857 => "11111111111110111111110111111000",
10858 => "11100011111101101111111011110101",
10859 => "11111000111111011111101011111011",
10860 => "11111101111111001111011011110111",
10861 => "11111000111111101111001100000000",
10862 => "11111110111101101110100111111000",
10863 => "11111010111101111111101111111111",
10864 => "11110010111010011110110111110100",
10865 => "11111100111101100000010011110101",
10866 => "11101110111101101111011111111011",
10867 => "11110010111010001111011111111100",
10868 => "11100010111110001111111011111011",
10869 => "11111000111011111111011011111011",
10870 => "11101011111101001110001011110101",
10871 => "11111011111110011111010111111110",
10872 => "11101100111000010000010100000000",
10873 => "00000000111010110000010011110111",
10874 => "11101010111100101111011111110110",
10875 => "11110010111000001111010111111111",
10876 => "11100000111010001111110000000001",
10877 => "11111101111001111111000011111010",
10878 => "11101010111100011111001011110111",
10879 => "11110001111110011110110011111010",
10880 => "11100110111111011111010111111000",
10881 => "00000001111000100000000111110101",
10882 => "11101001111101011111100111110101",
10883 => "11110111111010101111001100000000",
10884 => "11100001110111001111100011111010",
10885 => "11110101111001011110010011110001",
10886 => "11101100111100011110110111111001",
10887 => "11110100111110111110110111111100",
10888 => "11110001000001101110010111110010",
10889 => "11111101111011001111111011110101",
10890 => "11111010111101111111010111110100",
10891 => "11111011111110111111011111111110",
10892 => "11110111111001101111010111110110",
10893 => "11101110111010011111011111110111",
10894 => "11101111111010011111011111110011",
10895 => "11111010111101101110110111111011",
10896 => "11101000111111011111000111110001",
10897 => "11111101111001110000010011110010",
10898 => "11111000111110011111101111111101",
10899 => "11111010111010011111011100000010",
10900 => "11110001111001101111001011111010",
10901 => "11110000111010111111110111111110",
10902 => "11111000111110101111011011110110",
10903 => "11110010111110101111011011111011",
10904 => "11111100111101011111100111110010",
10905 => "11111100111111001111110011110110",
10906 => "11110110111100011111010111110011",
10907 => "11110101111101101111110000000010",
10908 => "00000110111101011111001111110101",
10909 => "11110100111110011111010000000000",
10910 => "11111001111101101111100011111001",
10911 => "11110110111111101111000111111001",
10912 => "11101111111010001111100011110011",
10913 => "00000000111101011111111011111101",
10914 => "11111001111111011111011111111001",
10915 => "11101110111010110000000000000000",
10916 => "11101000111011101110110011101001",
10917 => "11101110000000001111100111111100",
10918 => "11101001111111111110011111111001",
10919 => "11111111111110111111000111111001",
10920 => "11110111111001000000010100000111",
10921 => "11111011111101100000000011111100",
10922 => "11101111000000101111100011111010",
10923 => "11110110111111111111101000000001",
10924 => "11111000111001101111110100000110",
10925 => "11111011111101001111101011110101",
10926 => "11101011111111001111100011110101",
10927 => "00000000000000001111001011111010",
10928 => "00000011000000100000001100000100",
10929 => "00000010111110001111111111111101",
10930 => "11011100111100111111101011101011",
10931 => "11110111111110101111111100000011",
10932 => "11111000111110010000011000000011",
10933 => "00000110000000001110111111111011",
10934 => "00000010111111000000100111110111",
10935 => "11111110111111001111110011111100",
10936 => "00000100111011101111110111111011",
10937 => "00000001000000100000001000000000",
10938 => "11101001111101011111101011110001",
10939 => "11111000111111101111110011111101",
10940 => "11111111111011111111010111111011",
10941 => "11101011000000111111100111111010",
10942 => "11111101000000001111000011110101",
10943 => "11111110111111011111110011111111",
10944 => "00000001111110011111110111111100",
10945 => "11110111000000011111110100000000",
10946 => "11110001111110011111011111110101",
10947 => "11110101000000011111101111111111",
10948 => "11111001111111001111111011111100",
10949 => "11111011111110001111101111111100",
10950 => "11111100111111101110110111111000",
10951 => "11111100111110101111111111111000",
10952 => "00000000111101010000001111111000",
10953 => "11110110111111111111111011111000",
10954 => "11110001111110111111101011111001",
10955 => "11111000000000011111100011111010",
10956 => "11111010111101001111111111111100",
10957 => "00000000111010000000010011110110",
10958 => "11111000111100001110001011110111",
10959 => "11110011111110001111111011110110",
10960 => "11111111000001011111111100000101",
10961 => "11100100000010000000000111111010",
10962 => "00000111111111011111101000000101",
10963 => "11111001111111100000000111111000",
10964 => "11111101111011101111101100000011",
10965 => "00000001000010110000010011110000",
10966 => "11111000000001101111111011111000",
10967 => "00000001000010101111100111100000",
10968 => "11101111111100111111111100000111",
10969 => "11010001111110111111011100001001",
10970 => "00000010111111011101111111111101",
10971 => "11110111111010101111111011100110",
10972 => "00000010111001101111110111110111",
10973 => "11111011111111111111100111001110",
10974 => "00000000000001000000011011111001",
10975 => "00000100000000101111110011010110",
10976 => "11101101111011111111101111111111",
10977 => "00000111111010010000100000000000",
10978 => "11110111111110100000100111110100",
10979 => "11110011111111101111100011101100",
10980 => "11110010111001101111011100000000",
10981 => "11110111111100111111001011110101",
10982 => "11111001111110011111111111111001",
10983 => "11111110111110001111100100000010",
10984 => "11110110000000110000100000001010",
10985 => "00010000000001110001001111110001",
10986 => "00000000111111100001100000001001",
10987 => "11110011000001011111100100000001",
10988 => "11111011111100100000001100010010",
10989 => "00000000111111000000001100010010",
10990 => "00000101000001110000000011110110",
10991 => "11110111000010101111111100010111",
10992 => "11110111000000010000001100000111",
10993 => "00001110000000100000000111111001",
10994 => "11111101111110010000111100000011",
10995 => "11110111000000001111111100000011",
10996 => "11111011111100001111101111111110",
10997 => "11111011000001010000010000000011",
10998 => "11111111111111100000001011111000",
10999 => "00000011000000010000001100010011",
11000 => "11110101000000011111101000000011",
11001 => "11111010111110001111011111111111",
11002 => "00000011111111111111011000000110",
11003 => "11110110111110010000001111111110",
11004 => "11110101111110100000000111111011",
11005 => "00000010111111110000000011111011",
11006 => "11110110000000011111111111110101",
11007 => "00000110000000011111101011111001",
11008 => "11110010000001111111111100000100",
11009 => "00000110111001101111110111111000",
11010 => "00000011000000110000101011111100",
11011 => "11111110111110011111010011111111",
11012 => "11110110000011100000000000000001",
11013 => "00000011111101011111000100001011",
11014 => "00000110111111100000000011110101",
11015 => "11111010111110101111100100001010",
11016 => "11101011111110011111010100000010",
11017 => "00011010111100000000100111111111",
11018 => "00001110111101110001011100001001",
11019 => "11111011111101011111001000000001",
11020 => "11111111000001011111100100000101",
11021 => "11111010111111100000011100001110",
11022 => "11110100111101110000010011110011",
11023 => "11111001111110111111000100010010",
11024 => "00000100111111011111100000000011",
11025 => "00001100000000010000000011111000",
11026 => "11110011111110000000110111101101",
11027 => "11111101000000111111111100000000",
11028 => "11111010111101010000000011111010",
11029 => "11111110111101001111111000001101",
11030 => "00001001111110010000001111111000",
11031 => "11111011111111010000001100001010",
11032 => "00001011111101101111010011111000",
11033 => "11110110000011001111100111111001",
11034 => "00000101111100001111110100000000",
11035 => "11110010000010010000101100000011",
11036 => "11111011111110101110111111101100",
11037 => "11101001111110010001001100000101",
11038 => "11111000000011001111100111111001",
11039 => "11111111111111101111010100000001",
11040 => "11111111000000101111100111110001",
11041 => "11110010111111101111001111111100",
11042 => "00001001111100101111110100000101",
11043 => "11110100111100101111111100000000",
11044 => "00000011111110111111110011111001",
11045 => "11111110111111011111110111111101",
11046 => "11110110111111011111101111110011",
11047 => "11111011111111101111011000000110",
11048 => "11110101111110101111110011110101",
11049 => "11110110111110001111110011110110",
11050 => "11101101111110011111010011110011",
11051 => "11110100111110101111101100000010",
11052 => "11111010111110011111101011111111",
11053 => "11110110111011111111000111111001",
11054 => "11111001111110101110101011110111",
11055 => "11111010111111001111111011110010",
11056 => "11110011111101101111101100001100",
11057 => "11010000111110100000001000000011",
11058 => "11110101000000101100010011111010",
11059 => "11111000111110111111110111110101",
11060 => "00001010111011010000001111111100",
11061 => "11111101111111010000101111101001",
11062 => "11111101000001110001001111110010",
11063 => "11111111000000110000100011001100",
11064 => "11111000111011011111110000000100",
11065 => "11101001111010111110011000000101",
11066 => "00000110000001011101100000000101",
11067 => "11101111111110000000010011110101",
11068 => "11111101111000001111101000000010",
11069 => "11110110000000011111011111110101",
11070 => "11111011111111001111100011110110",
11071 => "00000001111111010000000011101000",
11072 => "11111101000010011111101100000100",
11073 => "00000001111111001111110000000111",
11074 => "00001001000001011111001100000111",
11075 => "11101111111111001111111111100101",
11076 => "00001000000011001111011100000100",
11077 => "11101100000010011111100011101101",
11078 => "00001010000000110000010111110000",
11079 => "11111111000000100000100011110111",
11080 => "11111001111110011111011100000110",
11081 => "00001000111011110000011000000001",
11082 => "11111111111110110000011111111001",
11083 => "11100011111111111111110111010111",
11084 => "11111011000110111111110000010001",
11085 => "11101000111110101111111111101111",
11086 => "11111000000000100000101111110010",
11087 => "11111011000000001111100011111111",
11088 => "00000101111001100000011000001010",
11089 => "00001010000000110000100111111101",
11090 => "11111111000011010000111111111111",
11091 => "11101000000001000000011100001100",
11092 => "00000000111110101111111000001010",
11093 => "11111101000000110000110000000100",
11094 => "11111001000000110000101011100011",
11095 => "00000100000000010000010100001011",
11096 => "00001100111101010000010000000100",
11097 => "00010001000010000000100011111110",
11098 => "11110101000100110001011111111100",
11099 => "11101110000010100000001011110101",
11100 => "11111000000010101111101100001101",
11101 => "11110010111111111111111000001100",
11102 => "11110011111111010000101011100001",
11103 => "00000110111110000000011100001000",
11104 => "00001000111111101111111111111110",
11105 => "00001010000000101111111000000010",
11106 => "11111110000010110000101111111011",
11107 => "11110111000010100000000111100111",
11108 => "00000001000000010000001100010010",
11109 => "11111010111110110000011000001010",
11110 => "11110001000000110000101011010111",
11111 => "11111110000010010000100100000001",
11112 => "00000010000001010000011100000010",
11113 => "00000001000100001111010111111101",
11114 => "00001011000010100000011000000101",
11115 => "11110011000011010000010111111110",
11116 => "00001011000000011111110100010000",
11117 => "00000101000001000000111000001110",
11118 => "00001100000010010000011111010101",
11119 => "00001001111111011111101100000011",
11120 => "11111001000010001111111100000110",
11121 => "11111110000000001111100100000010",
11122 => "00001100000011100001001000000001",
11123 => "00000101111111101111111000100000",
11124 => "11111001000010000000011100000110",
11125 => "00000111000011011111100000001010",
11126 => "11110110111101100000101011110011",
11127 => "00001001111110101111010000001111",
11128 => "00000001000000011111101000001010",
11129 => "00001100000001100000101011111111",
11130 => "00000111000001000001001000000000",
11131 => "11111010111101011111111100001011",
11132 => "11111110111110000000101111111111",
11133 => "00001011111111110000111100011001",
11134 => "11111011111111110000100011101010",
11135 => "00000110000000001111111100010001",
11136 => "11111001000000001110110000001000",
11137 => "00000110000000010000011000000110",
11138 => "00000101000001101111111100000000",
11139 => "00000001111110011111101011111101",
11140 => "11110111000000010000010000000001",
11141 => "00000011000011111111100011110111",
11142 => "11111010111110010000110011110011",
11143 => "11111101000000011111011011111111",
11144 => "00000100000000101111011011111011",
11145 => "00001010111100110000001000000001",
11146 => "11110100000100010001000111110010",
11147 => "11101111111111111111101111111001",
11148 => "00001100000000011111010111110111",
11149 => "11111010000001100001001000001110",
11150 => "00001011111111111111011011110111",
11151 => "11110101111111000000111000000110",
11152 => "00000100111011011111100011111101",
11153 => "11100011000000111111101111110110",
11154 => "11111111111101001101100111111101",
11155 => "11110100000000101111110000000001",
11156 => "11110010111010101111011011111101",
11157 => "11101101111111110000000000000011",
11158 => "11110000111111011110010111110111",
11159 => "11111001111111101111101111101101",
11160 => "00001110111011110000100100000001",
11161 => "11111010000010001111011111111110",
11162 => "11111101000000111111100111111011",
11163 => "11110111000001100000001111111000",
11164 => "00001101111100101111011111110101",
11165 => "00000000111110100000111111111100",
11166 => "00000010000000100000001111110101",
11167 => "00000011000000011111111011111110",
11168 => "11111101111110111111111000000110",
11169 => "00001111000100011111010000000100",
11170 => "00001001000011100000011100001010",
11171 => "11101110000000101111111011110010",
11172 => "00000111000000001111010100000001",
11173 => "11110110000010000000101111110110",
11174 => "00000011000011010000001111110011",
11175 => "00000101000000101111110100001001",
11176 => "00000100000010010000001000000100",
11177 => "00010110000000000000001000000011",
11178 => "00001101000001100001010000001100",
11179 => "11110110000010011111111111110010",
11180 => "11111100000000101111011100001100",
11181 => "11110000000000011111111000000100",
11182 => "00001100000001110000100111110010",
11183 => "00000000000000011111111100011101",
11184 => "00001111111111000000101111111100",
11185 => "00000110000100111111100000001000",
11186 => "00001001111111000000001000000011",
11187 => "11101101000101010000011111100011",
11188 => "11111011111111101111101100010101",
11189 => "11110110111111100001000011111110",
11190 => "11111010000011010000101011100111",
11191 => "00000100111111100000110000000101",
11192 => "00010011111011010000010111111010",
11193 => "00000110000100001111011100000011",
11194 => "11111010000000000000011011111100",
11195 => "11101000000010100000010111110001",
11196 => "00000100111100110000001000000011",
11197 => "11111110111110100001011100001000",
11198 => "00000011000011100000110111010010",
11199 => "00000000111110110000001000000010",
11200 => "00000011111111010000001111111001",
11201 => "11111100000001111111110111111010",
11202 => "11110011000000100000000111110100",
11203 => "11100111000010111111110011110001",
11204 => "00000010000001010000011100001010",
11205 => "00001110111110010000100011111100",
11206 => "00000010000011000000010110110001",
11207 => "11111011000000110000001111110100",
11208 => "00001001000000110000011111111010",
11209 => "00000010000100001111001000000100",
11210 => "11110101000001100000100111111111",
11211 => "11101000000011000000000000000110",
11212 => "00000110111111010000000100000101",
11213 => "00000110000000100001000000010001",
11214 => "00001111000000110000010010011101",
11215 => "00000000000010000000101000000000",
11216 => "00000011000001010000010111111100",
11217 => "00000000000001111110100100000011",
11218 => "11111101000000100000010111110111",
11219 => "11111111000000111111110100000010",
11220 => "00000101111111001111110000000111",
11221 => "00001101111111010000110000001100",
11222 => "11111111111110000000001011000110",
11223 => "00000000111111111111111000000100",
11224 => "11111010000001110000010011111111",
11225 => "11111011000010101111010100000101",
11226 => "11111001000000010000010111111100",
11227 => "00000101000000001111111100000110",
11228 => "00000110000001110000010111111101",
11229 => "00001100111111100000111000000000",
11230 => "00000100111110110000111011001110",
11231 => "00000010111111110000011100000101",
11232 => "11111100000000011111111111111111",
11233 => "11111011000001111111101100000001",
11234 => "00000110000000111111100000000010",
11235 => "00001111111110100000010100010001",
11236 => "00000101111111100000011100000000",
11237 => "00001010000001000000011011111101",
11238 => "00000111000000100000111011110011",
11239 => "00000010111110001111110100000000",
11240 => "00000001000010011111110000000000",
11241 => "11111110000100010000000000000010",
11242 => "11111111000001010000001111111010",
11243 => "11110101111110010000011000000000",
11244 => "00000011000001000000010100000110",
11245 => "00000101000011010001000100000010",
11246 => "11111111000010100000010011110010",
11247 => "00000000000001111111101111111110",
11248 => "11111001000001011111100011111110",
11249 => "11110000111100101111000111111010",
11250 => "11111001111111011111001011111000",
11251 => "11111010111100001111110111111010",
11252 => "00001011111111101111110011111110",
11253 => "00000001000000101111010111101111",
11254 => "00001110111101010000001011111000",
11255 => "11111110111111111111111011111000",
11256 => "11110001111110001111100111111010",
11257 => "11111110111100000000000011110110",
11258 => "00000100111101101111100000000000",
11259 => "11111000111110001111010111111101",
11260 => "11110101111011000000000100000100",
11261 => "11110001111111001110101111111111",
11262 => "11101111111110101110000011110101",
11263 => "11110110111111101111110011111100",
11264 => "00000111111010000000001111111001",
11265 => "11111100000001001111011011111101",
11266 => "11110010000001000000001111111010",
11267 => "11111000000000010000001011101110",
11268 => "00001000111001011111101111110100",
11269 => "11110001111100010000101111110111",
11270 => "11111011111111110000010111110101",
11271 => "00000111111111010000011011111100",
11272 => "00000111000111000000001011111110",
11273 => "11101111000011011110011000000101",
11274 => "00000100111111111111110000000100",
11275 => "11111011000000101111100011110101",
11276 => "00000110000101111110011000001000",
11277 => "11111011000001110000100100000001",
11278 => "00001001000000001111011111110010",
11279 => "11111101000000000000011011111110",
11280 => "11111111000011101111110100001000",
11281 => "11111011000100001110111000000011",
11282 => "00001000000000001111100100000000",
11283 => "11110101000010101111111011111100",
11284 => "00000110000101011111100000010111",
11285 => "11111011000000100000001100000001",
11286 => "00000100000001110001001111110000",
11287 => "00000011000001010000111011111001",
11288 => "00000101000100011111101100010001",
11289 => "11111110000011011110111000000011",
11290 => "00000001000000110000001100000000",
11291 => "11110000000000101111110011111111",
11292 => "11111110111111000000111011101110",
11293 => "00001010000000010000001100000000",
11294 => "00001001000001000001110011010010",
11295 => "11111110000001010000100111110111",
11296 => "00001110000101101111110100000011",
11297 => "11111010000110101110011100000101",
11298 => "11111101000000110001011011111101",
11299 => "00000101000001001111101100010011",
11300 => "00000001111111000001001111100111",
11301 => "00010100000001010001010100010101",
11302 => "00001000000011100000111110111010",
11303 => "11111101000001100000010011111011",
11304 => "00001011000010100000011011111010",
11305 => "11110110001000001110011111111100",
11306 => "11101100000001010000111011110111",
11307 => "11111011000010111111111000011010",
11308 => "00001110111100010001110011110001",
11309 => "00110001111101010010000100011001",
11310 => "00001111000100000001000011001110",
11311 => "11111110000001111111111000000101",
11312 => "11111101000101101111000000000001",
11313 => "00000001000011001111010000000000",
11314 => "11110111000010010000100000000000",
11315 => "11110011000010001111101100001000",
11316 => "11111101000000100001101100000010",
11317 => "00101010111110010000011100010001",
11318 => "00010100111111100010001110110101",
11319 => "11110101000000101111111111111010",
11320 => "00000101111111110000000111111100",
11321 => "00000101000001100000110000000100",
11322 => "11111001000000100001000000001010",
11323 => "11001010000000111111100111110100",
11324 => "11111110000001011110110100001010",
11325 => "11111101111111000000100100000110",
11326 => "11111101111111110001011011000100",
11327 => "11111000000001011111111100000001",
11328 => "00000101000000000000100100000100",
11329 => "00001001111111100000110100000100",
11330 => "00010001000010000001001100001111",
11331 => "11101011111111010000000000001011",
11332 => "00000100000001110000010000001101",
11333 => "00001000000010100001001000000011",
11334 => "00000001000010110001010111011001",
11335 => "00000011000000110000010000001000",
11336 => "00000001000001010000101111111001",
11337 => "00001100000000110000001111111010",
11338 => "00010110000100110000100000001000",
11339 => "11111101000011010000100100001001",
11340 => "00001000000000000000100100011000",
11341 => "00000110000001000000100000001111",
11342 => "11111111000001100000011011101000",
11343 => "00000001000001101111111100001111",
11344 => "00000110000001000000110100000001",
11345 => "00000100000110110000010000000010",
11346 => "11111110000010111111110000000000",
11347 => "11110111000100110000101000000100",
11348 => "00001000000000011111110011110101",
11349 => "00000101000001100000111011111111",
11350 => "00000010000011000001001011110100",
11351 => "00000111000001010000101100000000",
11352 => "00000000000101000000100011110110",
11353 => "00001000000000110000001011111011",
11354 => "11110100000000110000100011101111",
11355 => "00000010111111000000000100001010",
11356 => "00001000000010110000001111111100",
11357 => "00010111111111100000011100001001",
11358 => "00001001000000010000001111111000",
11359 => "00000111111110100000001000001001",
11360 => "00000110111110111111100000000011",
11361 => "11100100000010000000000111111110",
11362 => "11111110111111001110110100000100",
11363 => "11110110111111111111110100000100",
11364 => "11111000111101101111011100000101",
11365 => "11110110000000000000001000000010",
11366 => "11110110000000101110011111110011",
11367 => "11111111000000001111011011101101",
11368 => "00000101111001000000101111111100",
11369 => "11111100000011101110101011111111",
11370 => "00000010000001111111110111111101",
11371 => "11110000000010100000011100000001",
11372 => "00000101110111111111010111111111",
11373 => "11101100000000000000100000000101",
11374 => "11111100111111111111101111110100",
11375 => "00001010000000010000011000000101",
11376 => "00000101000110111111110100001000",
11377 => "00001000000100101110001000000111",
11378 => "00000001000001101111110100000101",
11379 => "11110011000000110000001000000110",
11380 => "00000101000000011110100011101001",
11381 => "00010000000011010000101100001101",
11382 => "00010011000001110000100011100110",
11383 => "00000111000010001111111000000111",
11384 => "00001000000010110000011000001010",
11385 => "11111000000111001101000000000010",
11386 => "11111110000010001111111111111011",
11387 => "11110100000100000000000100010011",
11388 => "11111101111100111111100011100010",
11389 => "00001100000001100001000100001110",
11390 => "00001100111110111111111111100010",
11391 => "00000010000010000000000111111111",
11392 => "00001111000101010000011011111000",
11393 => "11110100001000001100110000000101",
11394 => "11111011000001010000000111110110",
11395 => "00000100000100000000000000011010",
11396 => "00000111111111000000000011001101",
11397 => "00010010000010000001011000010001",
11398 => "00000100000001100000000011010100",
11399 => "11111111000000010000011111111001",
11400 => "00001111000101110000000111111100",
11401 => "11101010001011101100111100000100",
11402 => "11111101000010000000100011111000",
11403 => "00010110000100110000010000011111",
11404 => "00000001111011010000100111100001",
11405 => "00100001000001110010010000010010",
11406 => "00010001000110100000110011000001",
11407 => "00000100000100100000100111111010",
11408 => "00001011000011100000110111110011",
11409 => "11110001000110101100101111111111",
11410 => "00001001111111100000010011111010",
11411 => "00000111000001000000001000100111",
11412 => "00010000111010101111101011001011",
11413 => "00011100000011000010110100011111",
11414 => "00010001000010101111111011000110",
11415 => "00000010000011000000001011111101",
11416 => "00000101000010110000001111111100",
11417 => "11111001000100001111110100000111",
11418 => "00000101000001100000011000001010",
11419 => "11000011000000110000010011110010",
11420 => "00000111000010101111011000001001",
11421 => "00001011000000010001000111111001",
11422 => "00001111000100010001001011000011",
11423 => "00000000000001000000101111110111",
11424 => "11111001111110101111110000000010",
11425 => "00000110111111010001010000000011",
11426 => "00000011000000100000100111111110",
11427 => "11011110111110001111011011001001",
11428 => "11110101000010101111110100100110",
11429 => "11110110000000011111100011110000",
11430 => "11111011111111000001011011011101",
11431 => "11111101111111000000011111111100",
11432 => "11110101111101011111111000000000",
11433 => "00010010111010110001101100000001",
11434 => "00010010000010100000100000001100",
11435 => "11100010111111111111110011000111",
11436 => "11111011000010111111101000111000",
11437 => "11110000000000001110100111101110",
11438 => "00001100111011010000101011101001",
11439 => "11111111111111010000100011111011",
11440 => "00000111111111110000101100000000",
11441 => "00001110000001010001010000000100",
11442 => "00100001000011100001010000010110",
11443 => "11110100000010101111111111111001",
11444 => "00001001000010001111100100100010",
11445 => "11110100000101100000111100001100",
11446 => "00000010000100100001001111110001",
11447 => "11111100000101010000010100001100",
11448 => "00001000000001110000011111110100",
11449 => "11111111000011000000111100010011",
11450 => "11111011000000111111111100010000",
11451 => "11110011000000000001000111110010",
11452 => "00001000000011011111010011111101",
11453 => "11110110000010000000101011110111",
11454 => "00000010000011011111100011110000",
11455 => "00001000000011110000111111111000",
11456 => "11110110000100010000000111101101",
11457 => "00000000111110110000000100000110",
11458 => "11100111000001111111100011111001",
11459 => "11111000111111000000010000000100",
11460 => "00000000000100001111001111111101",
11461 => "00001111000000001111101111111011",
11462 => "00000010111111101101110111110010",
11463 => "00001100000000100000011011110111",
11464 => "11111110111110011111110011111101",
11465 => "00000011111111101111110100000010",
11466 => "00001000111111010000010100000010",
11467 => "11111010111110001111101000000100",
11468 => "11111011111110101111110111111100",
11469 => "11111001000001001110101100001010",
11470 => "11110111111111101110101011110011",
11471 => "11111001000000001111110000000101",
11472 => "00001111111001100000010011101111",
11473 => "11111100111101101111100111111100",
11474 => "11111111111100001111111011111110",
11475 => "11110111000000110000010111111100",
11476 => "11110011111101111110110111110010",
11477 => "11010110111111001111011011111111",
11478 => "00000000111111101101111111110101",
11479 => "11111011000000101111110011111001",
11480 => "11111111000110101111110111111101",
11481 => "00000101000000111111011100000000",
11482 => "11110010111100100000100111110110",
11483 => "00000011111101111111101000000101",
11484 => "00000101111110011111011111111101",
11485 => "00011111111101100000100000000111",
11486 => "00001011111111001111111111101111",
11487 => "11110111111111100000001100001011",
11488 => "00000000000011000000001000000010",
11489 => "11110010000011101101111111111111",
11490 => "11110100000000000000100011111110",
11491 => "11111110000001111111110000001111",
11492 => "11111000111101001111111111110011",
11493 => "00011000111101100000011000001001",
11494 => "11111111000000010000001111100101",
11495 => "00000011000001100000010011110111",
11496 => "00000111000100010000011111111101",
11497 => "11110110001000001100010000000101",
11498 => "11111011111111010000010111111110",
11499 => "11101101111111100000010100001110",
11500 => "00000100111101010000111111101001",
11501 => "00100010000001010001101000001001",
11502 => "00000111000100110001111011010101",
11503 => "00000101000011010000011011111110",
11504 => "00001010000100101111111111111010",
11505 => "11110011001000101101010000001010",
11506 => "00000000000011000000111011111101",
11507 => "00001110000101010000001000001011",
11508 => "00000100111100010000100011010011",
11509 => "00011100000001110001101100010010",
11510 => "00001010000001100000101111000011",
11511 => "00001001000010101111101100000000",
11512 => "00000010000101000000110111111010",
11513 => "11110011000101111101100100000010",
11514 => "11111000000010000000000111111000",
11515 => "11110001000000110000010011111110",
11516 => "00001101111110001111100111010001",
11517 => "00010111000000110001110100001111",
11518 => "00001100000101010000011011000101",
11519 => "00000100000010010001000000000111",
11520 => "00000001111110011111110000000101",
11521 => "00010011000001000000101000000110",
11522 => "00000000111111000000101011111010",
11523 => "11000100000001011111111111011111",
11524 => "11111010000001011111000000010100",
11525 => "11110001111111101111110011111110",
11526 => "00000111111111010001000011000000",
11527 => "11111101000000110000111000001000",
11528 => "00001000111110011111100000000000",
11529 => "00010011000011010001100000000100",
11530 => "11101011111111110001111111110000",
11531 => "11101000000011100000001011110101",
11532 => "00000000000010101111111100101101",
11533 => "11111000111101010000100000010001",
11534 => "11111011000001010001000111011100",
11535 => "00000100000000100000011100010100",
11536 => "00001000111100111111111011111111",
11537 => "00001001000010010000111000000101",
11538 => "11100101111101100001000011101001",
11539 => "11110011000000111111110011101010",
11540 => "11110111111111000000110100011000",
11541 => "00000010111111001111101000000100",
11542 => "11111001111111010001101011101110",
11543 => "11111101111110101111110100000110",
11544 => "11111100111100110000000011111001",
11545 => "00001000000010100000110000000110",
11546 => "11101101111110110001011111110100",
11547 => "11111101000001110000000111111010",
11548 => "00000000000000100000101011111110",
11549 => "11110000000001100000000100001010",
11550 => "11110101111111100001000111111000",
11551 => "11111010111111010000000111111111",
11552 => "00000100111101100000110111101100",
11553 => "00000111000000010000010011111111",
11554 => "11111100111110000000100111110010",
11555 => "00000010111111100000100011101111",
11556 => "00000001111101101111101111111101",
11557 => "11101011111110010000000111111111",
11558 => "11111000000000101111110111111000",
11559 => "00000000111111101111111000000010",
11560 => "00000100000000011111011011101011",
11561 => "11110110111110111111101011111010",
11562 => "11100100110101011111010011101111",
11563 => "11110101111100000000000111101100",
11564 => "11111111111111111110111000001111",
11565 => "11101010111111011110110111101111",
11566 => "00000000111100011111001011110101",
11567 => "11111010111101110000010111110111",
11568 => "11111000111111101111100011111101",
11569 => "00000001000000011111111011111011",
11570 => "11110101111110111111110011110111",
11571 => "11110101111111101111110100000001",
11572 => "11110111111110101111011111111011",
11573 => "11110111111101101111101111111101",
11574 => "11111101111100111111000011110011",
11575 => "11111101111110101111100111111011",
11576 => "11101100000000001111110011111010",
11577 => "00000100111011001111011111110110",
11578 => "00000101111101011111100011111111",
11579 => "11111101111011101111000100000101",
11580 => "11110000111110011111100011111000",
11581 => "00000101111111101111010100000001",
11582 => "11111100111100011111000111111001",
11583 => "11110011111011111111011100000001",
11584 => "00000101111101011111111100000110",
11585 => "11111111000100011111001100000001",
11586 => "00000010111111101111101100000011",
11587 => "11110011000011010000011111110010",
11588 => "00000001111010111111010100001011",
11589 => "11011010111111000000100011111000",
11590 => "00001000000100000000100111110010",
11591 => "00000011000001100000011011111110",
11592 => "00000101111110101111101100000111",
11593 => "11111100000001101111110000001111",
11594 => "00001001111110000000001100001101",
11595 => "11110101000000011111110111111000",
11596 => "00000100000001101111011000000010",
11597 => "11101001000001010000000100000000",
11598 => "11111100000011010001001011100110",
11599 => "11111110000010000000011011111010",
11600 => "00000110000101110000000000000111",
11601 => "11111111000010011111001100001000",
11602 => "00000111000010000000011100001011",
11603 => "11000110000001010000010111110010",
11604 => "00000011000001011110110111111110",
11605 => "11110000000001010001001000000110",
11606 => "00001001000010000000100011011100",
11607 => "00000011000011110000000011111011",
11608 => "00000100001010001111011100001101",
11609 => "11111011000100011111010100001011",
11610 => "00010010111111010000011000001110",
11611 => "11100011000000000000011011100010",
11612 => "11111110000100011111110111111111",
11613 => "00001001000011000000111000001001",
11614 => "00001000000010010001101010110111",
11615 => "00001001000010011111111111111001",
11616 => "00000111000000000000010100001010",
11617 => "11111010000010011111001100001101",
11618 => "11111010000000101111101000000000",
11619 => "11001000000000100000001111100010",
11620 => "00001101000001101111001011101110",
11621 => "11111100111111000001001000000100",
11622 => "00001111000000010001000011001111",
11623 => "00000110000000100000110111111010",
11624 => "00000110111111010000010000000100",
11625 => "00000100000100111110111011111111",
11626 => "11100010000000110000101111101011",
11627 => "11110111000001111111110111111111",
11628 => "11110000111111100000101100000001",
11629 => "00010001111101110000110000001010",
11630 => "11110101000011000000110011001000",
11631 => "00000000000000100000000000000001",
11632 => "00000000111111111111100111111000",
11633 => "00001000000000100000011011111111",
11634 => "11101110000000100010000011101010",
11635 => "00001101111110111111110100001001",
11636 => "11111110111111000001001111110101",
11637 => "00010101111110000000001100010001",
11638 => "11111101000000010001100011100101",
11639 => "11111100111110100000000100010001",
11640 => "11111101111110011111110011100100",
11641 => "11111111000010011111010111110010",
11642 => "11010111111111110000111111011110",
11643 => "00001000000000011111100100000101",
11644 => "11111111111011110000100111101010",
11645 => "00001100111011100000100100001010",
11646 => "11110110000000000000000011110011",
11647 => "11111000111110011111111000000110",
11648 => "11111101111011111111110111101111",
11649 => "00001000000010110000000111110001",
11650 => "11111111111101000001110111111011",
11651 => "00000101000010011111101100010100",
11652 => "11111001111010110001000111101001",
11653 => "00000010000011010000110100011000",
11654 => "11101110000000000000010111111011",
11655 => "11111001111111001111001000001111",
11656 => "00000101111101010000001111110110",
11657 => "11100110000011111110110111111110",
11658 => "00000111111111001111011000000010",
11659 => "11110111111111000000001011111111",
11660 => "11111101111011011111110111101101",
11661 => "11111010000001010001011100000100",
11662 => "11111010000011000000010011111000",
11663 => "11111011000010011111100011110011",
11664 => "11110111000001100000000011110010",
11665 => "11101101111010001111001011111110",
11666 => "11101001111010001101111011110111",
11667 => "11111000111010011111100011110101",
11668 => "00000100000000011111010111101001",
11669 => "00000110111100011111110111101100",
11670 => "00001010111110010000000011110101",
11671 => "11111101111111010000001011100010",
11672 => "11101111111111111111101111101001",
11673 => "11111000111000100000000111110011",
11674 => "11011111111011011111001011100100",
11675 => "11111001111011001111011111111010",
11676 => "11110111111111011111011011110011",
11677 => "11110111110111011110110011110101",
11678 => "11111010111010101110110011110110",
11679 => "11110000111010011111011011110101",
11680 => "11110101000000100000000100001001",
11681 => "11110000111101101111110011110101",
11682 => "00000000111110101111011111111011",
11683 => "11111101111101001111100111111011",
11684 => "11111010111111101111100000000001",
11685 => "11010010000010001111101111111001",
11686 => "11111000000001001111011111110111",
11687 => "00000001000000011111100111110010",
11688 => "11110100000000011111101000000100",
11689 => "00000000111111110000000000000110",
11690 => "00001100000000001111001100001111",
11691 => "11101011111101101111011111101011",
11692 => "00000101111110101110100100000110",
11693 => "11010101111111111111010111110111",
11694 => "00010100111110110000000011110001",
11695 => "11111101111111000000110011111000",
11696 => "11111111000000011111011000010000",
11697 => "00000001111110100001000100001010",
11698 => "00010100000000001111010100001101",
11699 => "11010000000000111111100111011100",
11700 => "00000001000110001110010100010101",
11701 => "11000110000000000000001011111000",
11702 => "00000111000001110000111111100101",
11703 => "11111110000010010000110011101100",
11704 => "11111110000101100000000000001010",
11705 => "00000001111111110000011100001111",
11706 => "00001110000001101111000100010111",
11707 => "10111000111111010000001111011000",
11708 => "00001111001000011100110100010010",
11709 => "11001100000010110001001011111011",
11710 => "00001001000001010000001011001110",
11711 => "00000000000010100000111111110010",
11712 => "00001010000100110000000100001011",
11713 => "00000101000011101111100000001001",
11714 => "00010111000010111111100100010111",
11715 => "10101100000001100000011111100011",
11716 => "00001101001000001100100000000111",
11717 => "11011001000011010001000100000111",
11718 => "00000110000001100000101111000000",
11719 => "00000110000001100000110011110101",
11720 => "00000111000011110000001011111101",
11721 => "00000011000010101110111111111111",
11722 => "11110100000010101111001011111010",
11723 => "11001100000001000000001111100111",
11724 => "00001000000100001110101111110111",
11725 => "00001011111111000001011100000101",
11726 => "00001111000011101111000110111100",
11727 => "00000001000000110000001111111001",
11728 => "00000101000000011111101111111001",
11729 => "11111010000100001110000100000010",
11730 => "11111100000001100000110111110111",
11731 => "00010000000000101111011000010110",
11732 => "11111000111100000000110111101001",
11733 => "00010101111111100001001000010000",
11734 => "11111110000000100000101011010110",
11735 => "11111001111111101111101100001000",
11736 => "00000010000010101111101111101111",
11737 => "11111011000010101111010011111000",
11738 => "00000000111110100001000111111001",
11739 => "00010001000001101111110100010100",
11740 => "00000000000000010001011111101010",
11741 => "00011110111111010001001100001010",
11742 => "00000000111111110000100011101000",
11743 => "11111010111100101111011100000110",
11744 => "00000100000001111111111111110101",
11745 => "11110001000001101110001011111101",
11746 => "00000001111101010000010000000100",
11747 => "00001010111100111111010100010010",
11748 => "11111101111101000001000111100001",
11749 => "00011100111111100001010000000101",
11750 => "11111011000010000000110011111000",
11751 => "11110110000001101111011111111111",
11752 => "11111100000000010000000011110101",
11753 => "11100111000000101100110100000000",
11754 => "00001011111101011110000100001001",
11755 => "11111111111110101111110011111010",
11756 => "11111011111011100000011011101010",
11757 => "00001101000011000000011111111001",
11758 => "11110110000000100000010011110100",
11759 => "11111000000011101111110011101000",
11760 => "00000001000000100000001011111001",
11761 => "11101011000001101110100100001001",
11762 => "00000011111110011101111000010100",
11763 => "11110101000000011111101011100110",
11764 => "00001110111110101111011111011000",
11765 => "00000110000010000001001011100100",
11766 => "00000011000010101111111111110010",
11767 => "11111010000100100000100111010110",
11768 => "00000000000011001111011111110010",
11769 => "11111011111110110000000111110111",
11770 => "11101101110111001111000111110111",
11771 => "11110110111100010000000011111111",
11772 => "11111000000100011111011111110100",
11773 => "11111110111101011101101111101010",
11774 => "11111111111011101111010111111000",
11775 => "00000011111110001111101111101110",
11776 => "11101101111111011111010011101011",
11777 => "11101001111001101111110011110101",
11778 => "11100101111100001101110011101000",
11779 => "11110011111011111110111111101110",
11780 => "11111011111101001111110011110100",
11781 => "11111001111001101110110011101001",
11782 => "11111010111001111110110111110110",
11783 => "11110000111010101111001111101100",
11784 => "11110110111001010000000011111110",
11785 => "11100110111011001110001011111101",
11786 => "00000011111111111110101111111101",
11787 => "11110111111111101111101111111001",
11788 => "11111101111001011110111011110100",
11789 => "11010000000000001111001111111100",
11790 => "11110011111101101111100011110100",
11791 => "11111011111111010000000011110001",
11792 => "11111111000101110000011100000111",
11793 => "11110001000001111101101100001001",
11794 => "00001000000001011110100000001001",
11795 => "11101000000000011111111011101101",
11796 => "00000011000000111110011000000011",
11797 => "11101110000001110000100111110101",
11798 => "00001011000010100000000111101111",
11799 => "00000101000010000000001111110100",
11800 => "00000111000111000000000100001011",
11801 => "11110011000000011111000000001101",
11802 => "00001011000000001110100000001000",
11803 => "11011101111111000000001011100010",
11804 => "11111110000110111110101100000100",
11805 => "11101010000001111111110011110111",
11806 => "00000101000001010000111111100011",
11807 => "11111110000000110000000111110000",
11808 => "00001101001010000000000111111100",
11809 => "11110110000011011111010000000010",
11810 => "00000110000001111110110000001000",
11811 => "11001000000100000000001011101000",
11812 => "00000110001001011101110011110111",
11813 => "11110001000000000001010111111001",
11814 => "00001001000000100000011010111100",
11815 => "11111010000001010000011111100001",
11816 => "00001101000101110000101111111000",
11817 => "11101111000010011101100111111011",
11818 => "00001100000000001110101100010010",
11819 => "11010100000000100000000100001011",
11820 => "00010111000101011101111111111011",
11821 => "00000000000010010000110000010000",
11822 => "00011010000000011111101110101110",
11823 => "00000001000000100000011111110010",
11824 => "00000111000010000000011011110110",
11825 => "11110110000011111101100011111001",
11826 => "11111011000001100000000000000111",
11827 => "11010101000000101111111000010101",
11828 => "00001101000010011111001111111111",
11829 => "00001111111111000010000100010110",
11830 => "00001100000010001111001110110100",
11831 => "11111010000001010000000000000010",
11832 => "11111110000001101111110011111011",
11833 => "11111110000000101110111111111100",
11834 => "11111110000001100000011100000100",
11835 => "00000000000000011111001000000110",
11836 => "00001100000000000000000111101101",
11837 => "00100010111110000001010000010100",
11838 => "00001111000000011111110111011001",
11839 => "11110101111111001111101000000100",
11840 => "11111010000001101111100111111111",
11841 => "11110001111101111111001011111110",
11842 => "00000111111111111111010100001101",
11843 => "11110000111110001111010111110110",
11844 => "00001001000001001111100111101101",
11845 => "00000100000000000000101011111001",
11846 => "00001101111110010000010111011111",
11847 => "11110011000000111111111011111001",
11848 => "00000000000001001111101100000101",
11849 => "11110000111111001110010100001001",
11850 => "00001001111111001101111000010100",
11851 => "11110101111011111111110111100011",
11852 => "11111011111110101110111011110111",
11853 => "11111001000010000000010011100111",
11854 => "00000001111111110000011011101001",
11855 => "11111010000000111111111011100100",
11856 => "11111101000000110000000100000110",
11857 => "11111000111110101111010000000111",
11858 => "00010101000000001111000000001111",
11859 => "11110011000001111111100111110001",
11860 => "00000101000000011110111111101011",
11861 => "11111000000010110000001111111110",
11862 => "11111100111111100000100011101010",
11863 => "11111110000011110000001111110001",
11864 => "00001001000001000000000111110001",
11865 => "00000011111101011111111000001010",
11866 => "11110000000000010000010011111111",
11867 => "11110100000001011111110111101100",
11868 => "00001010000010001111001011111001",
11869 => "11110110111111110000011011111011",
11870 => "00001100000001101111110011110000",
11871 => "11110100000001010000011000000110",
11872 => "11110110111110011111010011111001",
11873 => "11111101111100101111111011111000",
11874 => "11101110111000011111001011110110",
11875 => "11110111111110101111110011111010",
11876 => "11101101111111001101100100001011",
11877 => "11101101111100111101011011110011",
11878 => "11101100111011011100011011111000",
11879 => "11111001111110011111100111101100",
11880 => "11110110111110001111110111100111",
11881 => "11100111111100110000000011110001",
11882 => "11100001111100001110100011100101",
11883 => "11110101111100011111001011110010",
11884 => "11110111111111001111010011111101",
11885 => "11111001111000111111000011101010",
11886 => "11111001111011101110010111111000",
11887 => "11111000111011101111100111101011",
11888 => "11111010111010110000000000001100",
11889 => "11110011111101111111011100000000",
11890 => "00000001111110001110110000000010",
11891 => "11110010111101011111111111110111",
11892 => "11111111110101001110110100000101",
11893 => "11011101000001001111011000000001",
11894 => "11111010000000000000100011110111",
11895 => "11111101000001111111101111110101",
11896 => "00000000000011011111110100000000",
11897 => "00000001000000111111010000001001",
11898 => "00001000000000111111111000000001",
11899 => "11101111000001010000011000001000",
11900 => "00000011111001101101001011100111",
11901 => "11110010000001000000100100001001",
11902 => "00000100000010010000000011101011",
11903 => "00000101000000110000100100000101",
11904 => "00000011000100111111111100000011",
11905 => "11111010111111101111000011111011",
11906 => "11111010000000011111101111111011",
11907 => "11101111000000010000100100000001",
11908 => "00000101111101111110100011011001",
11909 => "00001011000000001111110000000011",
11910 => "00001011000001101111101011101011",
11911 => "00000001111111001111011011111000",
11912 => "11111001000011011111110111110100",
11913 => "11110100000011011111001011111100",
11914 => "11111110000001001111110111111101",
11915 => "11110001111111000000000000010111",
11916 => "11111111000000111110101011011110",
11917 => "00010000000001000000011100001010",
11918 => "00000010000000001111100111001011",
11919 => "00000110000000100000000000000010",
11920 => "11111101000100100000010011110111",
11921 => "11111111000001011111000011110101",
11922 => "00000000000001110000110100000010",
11923 => "11110011111110101111110100100001",
11924 => "11111110000010001111011111110110",
11925 => "00010011000000000000101100010010",
11926 => "00010010111110000000011110110110",
11927 => "11111111111111101111110000000110",
11928 => "11111101000101000000001100000001",
11929 => "00001001111111011111110011111110",
11930 => "00001001000000100001000000001101",
11931 => "11011000111111011111101100010111",
11932 => "00000011000100101110111111111001",
11933 => "00001110000000110000101000000101",
11934 => "00001001111101110000100110111001",
11935 => "11111110000001001111101100000111",
11936 => "00000100000000100000000000000001",
11937 => "00000010000000000000100011111100",
11938 => "00010001000001001111111100001101",
11939 => "11000001000000101111111011101110",
11940 => "00000000000001001111110000001101",
11941 => "00000101000000000000110011111111",
11942 => "00001010000001110001010011011000",
11943 => "11111101000010101111111111111101",
11944 => "00000011111111110000011000000111",
11945 => "11111101111111111111111000000100",
11946 => "11111101111101111111100100001011",
11947 => "11100110111101101111101111100011",
11948 => "00000100111111101111100111110011",
11949 => "11111000111110110001000111111100",
11950 => "00000101000000000001010111100010",
11951 => "11111101111110011111110011110100",
11952 => "11111000111111110000011100001001",
11953 => "11111101111100101111011100000100",
11954 => "00001101111110111111100100001010",
11955 => "11101110111110010000000011101010",
11956 => "00000011111111011111000100001110",
11957 => "11110001111111010000000011110101",
11958 => "00001101000000000000000111110010",
11959 => "00000001000001110000000111111011",
11960 => "00000001000001000000010000001011",
11961 => "11110101111100111111111100001001",
11962 => "00001110111101111111110000001110",
11963 => "11101011111011101111101011011111",
11964 => "11111101000010011110110111111100",
11965 => "11110001000011001111111111110101",
11966 => "00000001111111111111100111101111",
11967 => "11111110000001010000011111111111",
11968 => "11110110000000111111101100000010",
11969 => "11110011111011001111100011111011",
11970 => "11110100111101011110111111100111",
11971 => "11110011111011111111011111110001",
11972 => "00000110000001111111011011110011",
11973 => "11111000111111101111001011101101",
11974 => "00010000111101101111100111110011",
11975 => "11111001111100011111111111110010",
11976 => "11110101111000101111000011110100",
11977 => "11101010111100001110110011111010",
11978 => "11101100111001011110000111110110",
11979 => "11111010110110101111011111111111",
11980 => "11110010111000101110110111110101",
11981 => "11011011111101001110111011101001",
11982 => "11101100111100001101011011110101",
11983 => "11110011111110011111011011101010",
11984 => "11111101111110101111100011111001",
11985 => "11110001111101111111011011110101",
11986 => "11110011111110101110111011110000",
11987 => "11111000111101111111011011101111",
11988 => "11111001111110011111011111111111",
11989 => "11111011111001001111011011101010",
11990 => "11111001111111001110110011111010",
11991 => "11111011111101011111101011101100",
11992 => "00000000111111001111101111110110",
11993 => "00000011111011111111110000000001",
11994 => "00000011111110101111110100000010",
11995 => "11111001111100011111110111111100",
11996 => "11111101110111111111001111100111",
11997 => "11110110000000011111101011111100",
11998 => "11111111111010111101111111110011",
11999 => "11110101111110100000000111111100",
12000 => "00001011000101110000100011110000",
12001 => "11111111000000010000000100000010",
12002 => "11110111111111110000011011111001",
12003 => "11110101000000000000011100001000",
12004 => "00001101111101111110011011100111",
12005 => "00000101000000100000100000001000",
12006 => "11111100000010001101001011111010",
12007 => "11111111000000001111100000000100",
12008 => "00000011111011010000010011110110",
12009 => "11111110000001111111100000000000",
12010 => "11111001111101100000001011110000",
12011 => "00000000111110111111111000000111",
12012 => "11111110111100001111111111010111",
12013 => "00101001000001000000101100001000",
12014 => "11111111000000001111100111110100",
12015 => "00000001111111011111100100000011",
12016 => "00000011111011100000011011101101",
12017 => "11111101000010011111011111111101",
12018 => "11110011111111100000001111101011",
12019 => "11111101000001000000010100000110",
12020 => "00000011111010000000001110100101",
12021 => "00101001111111010000101000000010",
12022 => "00000100000011001111111111110100",
12023 => "00000101111111111111100000000000",
12024 => "11110100111010011111110111110111",
12025 => "00001000111111101111101011111110",
12026 => "11111110111110000000011111101111",
12027 => "00001101111110111111110100000101",
12028 => "00001000111100100000011011100011",
12029 => "00011110000001100000101100001000",
12030 => "00000111000000000000001111011011",
12031 => "00000000000000000000010100000111",
12032 => "11111100111101100000001100000110",
12033 => "00001000000010100000000100000100",
12034 => "11101011000001100000000111100101",
12035 => "11101101000001010000000011110100",
12036 => "11111101111110100000010100000111",
12037 => "00000101000000011111110111111110",
12038 => "00000110000011000010001111100010",
12039 => "00000010000000010000000000000101",
12040 => "11111111000000000000001000001100",
12041 => "00000010111111010000010100000100",
12042 => "11111011000011000000000011111110",
12043 => "11100010000001011111111111101100",
12044 => "11111100000010010000010100100000",
12045 => "00000001000010001111011100000000",
12046 => "00001010000001000001111111011111",
12047 => "11111101000000110000010111111111",
12048 => "00000000111101010000001100001110",
12049 => "00000101111111001111111000000101",
12050 => "11110101000001110000000011110100",
12051 => "11011011111110110000000111110111",
12052 => "11110011000000011111111000001000",
12053 => "00000011000000111111001100000000",
12054 => "11111100111101100001000111100101",
12055 => "11111110000001011111111100001001",
12056 => "00001100111111010001000100001011",
12057 => "00001101000001100000101100000110",
12058 => "11101011000100100000101011110011",
12059 => "11100110000001110000100111111100",
12060 => "11111101000001111110011111110111",
12061 => "11110011000000110000010000001101",
12062 => "00001111000001101111110111110011",
12063 => "00000100000001000000100100010001",
12064 => "00000011111111100000011111111100",
12065 => "00001011111101000000001100000011",
12066 => "11101100000010100000001011110100",
12067 => "11110100000000100000010011111011",
12068 => "00000000000010111110101111110000",
12069 => "11110001111111011111011100000001",
12070 => "11111101111110101110011011110010",
12071 => "00001011111111100000011000000100",
12072 => "00000101000010101111011111111110",
12073 => "00001101000010010000001111110101",
12074 => "11101001111111110000010011101010",
12075 => "11110010000100110000001011101110",
12076 => "00000101000010011111010111111110",
12077 => "11111101111110010000001011111010",
12078 => "00001010111111011110101011110111",
12079 => "00000110111101101111111000000100",
12080 => "11110011111000001111001111110101",
12081 => "11100010111100011111001111111000",
12082 => "11101101111011011101111011111010",
12083 => "11110101111010011111100111111011",
12084 => "11110101110111101111110111110101",
12085 => "11100010111100001111001111100100",
12086 => "11101110111100001110010111110101",
12087 => "11110110111101001111101111101000",
12088 => "11111010111110111111100111111101",
12089 => "11110010111111001111110111111010",
12090 => "11101110111110111110101111111000",
12091 => "11110101111110001111110011111100",
12092 => "11111001111111011111100100000100",
12093 => "11111101111100001111110011111000",
12094 => "11111011111111011110110011110110",
12095 => "11111110111111001111110111110101",
12096 => "11110110111111111111000111110101",
12097 => "11101011111110001111010011101100",
12098 => "11110011111100101110111011110010",
12099 => "11110111111110001111100011110010",
12100 => "11110100111011011111100011111101",
12101 => "11111110111010001111010011110001",
12102 => "11110110111101011110001011111011",
12103 => "11110010111100111111011011101000",
12104 => "11111001111010011111011111101111",
12105 => "11110111000000011111010100000000",
12106 => "00000001111010111111001011111110",
12107 => "11111000111101001111100111110011",
12108 => "11110101111011001111101111110101",
12109 => "11111011111110111111110011111001",
12110 => "11111110111001011101011111110011",
12111 => "11111010111101011111100011110110",
12112 => "11111011110110001111110011101011",
12113 => "11110100111111111110111011111100",
12114 => "11100011111100101111011111101101",
12115 => "11111011111111111111111111111111",
12116 => "11111000111000010000001011100101",
12117 => "00000110111010110000001011111000",
12118 => "11101111111111101101111111110011",
12119 => "11111100111111101111101111110101",
12120 => "11111110110110110000001111101010",
12121 => "00000001000000011111110011111010",
12122 => "11101000111100100000000011101101",
12123 => "11111011111110011111101011111111",
12124 => "11111000111100100000010111101010",
12125 => "11111010111101000000000000000000",
12126 => "11111100111110110000000111111001",
12127 => "11111011111110011111111100000011",
12128 => "00000110110111000000101011101100",
12129 => "11111111111100100000000000000100",
12130 => "11011110111101100000001111100110",
12131 => "11110110000001010000010111111100",
12132 => "00000111111111011111001100000010",
12133 => "11011001111110010000101100000110",
12134 => "11110011000001011110100011111001",
12135 => "11111001000000010000000000000111",
12136 => "00000010111001110000001011101011",
12137 => "00000001111110011111111111110111",
12138 => "11010000111101010000001011101000",
12139 => "11111011000000000000000111110001",
12140 => "00000000000000001111001011111110",
12141 => "11010010111010110000010000000001",
12142 => "11111010000001111110100011110011",
12143 => "11111000000000101111110100000001",
12144 => "11111010111101011111101111100111",
12145 => "00000010000001001111110011111011",
12146 => "11110100111111111111110111111011",
12147 => "11110101000000110000011111110001",
12148 => "11110010000000001101111000000011",
12149 => "11000000000000100000010100000000",
12150 => "11111010000001111101001111110111",
12151 => "00000000111101001111010111111111",
12152 => "11101111111110111111001111110011",
12153 => "11111100000001111111111111111000",
12154 => "11010011111111001111110011101010",
12155 => "11110001000010011111111111110100",
12156 => "11110100111111101110111100000100",
12157 => "11101111111100001110101011110110",
12158 => "11110110111011101101101011110111",
12159 => "00000011111101001111111111111100",
12160 => "00010000111110000000110111110101",
12161 => "00001000111111110000010011111001",
12162 => "11100010111100010000101111100111",
12163 => "11111001000000101111111000000011",
12164 => "00000010000000011111100111110010",
12165 => "11111011111010100000011000000111",
12166 => "11111101000001001101000011110100",
12167 => "11111101000001100000100000000011",
12168 => "11111101111101000000000011110011",
12169 => "11111010111100000000001011110000",
12170 => "11100101111000010000010111101001",
12171 => "11111000111100101111101111111100",
12172 => "11111101111111111111111011111101",
12173 => "11010100110111101111110111111011",
12174 => "11111011111111011110011111111001",
12175 => "11110011111110011111110011111010",
12176 => "11111010111101111111100111110110",
12177 => "11110001111011001111101111111010",
12178 => "11110001111001101111110111110111",
12179 => "11111011111001101111101111111011",
12180 => "00000000111110101111100000000011",
12181 => "11011110111101010000000100000000",
12182 => "11110111000000101111001111110101",
12183 => "11101101111111101111100011111000",
12184 => "11111000111011111111100011111001",
12185 => "11101101111110011111011011111101",
12186 => "11111000111101011110011111111001",
12187 => "11110111111110001111100100000000",
12188 => "11111011111011001111100011111000",
12189 => "11110010000000011111100011110111",
12190 => "11111001111110101110110011111000",
12191 => "11110111111111111111100011110010",
12192 => "00000000000000000000000000000000",
12193 => "00000000000000000000000000000000",
12194 => "00000000000000000000000000000000",
12195 => "00000000111111100000000000000011",
12196 => "00000011111111100000010100000101",
12197 => "00001100000001000000000000000001",
12198 => "11111110000000001111111011111111",
12199 => "00000001111111110000000000000000",
12200 => "11111101000000001111111111111110",
12201 => "00000001000000010000101111111110",
12202 => "11111101000000110000000000000101",
12203 => "00000011000000111111111100000000",
12204 => "00000010111111010000011100000101",
12205 => "00001010000001000000000000000010",
12206 => "11111110000000101111110100000011",
12207 => "00000011111111110000000100000010",
12208 => "11111100111111100000001011111110",
12209 => "11111101111111000000111111111100",
12210 => "00000000000000010000000000000010",
12211 => "11111100000000010000001011111110",
12212 => "00000110111101110000011111111110",
12213 => "00000000000001101111111100000001",
12214 => "11111110111111001111110000000001",
12215 => "00000100111111000000001000000011",
12216 => "00000000111110001111110111111101",
12217 => "11111111111111000000110100000000",
12218 => "11111001111101100000000100000010",
12219 => "11111111111110100000000011110111",
12220 => "00000100111111110000010000000000",
12221 => "11111110111101000000001111111001",
12222 => "11111110111111111111111000000011",
12223 => "11110101111101001111111000000010",
12224 => "11110101111111011111001100000010",
12225 => "11111000111111010000100011111110",
12226 => "11111111111110101111101011111111",
12227 => "11110111111110011111011111110001",
12228 => "11111110111111100000011111110101",
12229 => "11100001111101101111100111110110",
12230 => "11111111111101011111010111111101",
12231 => "11111101111100101111100111111010",
12232 => "11100111111100101111010011111111",
12233 => "11111001111101101111110011111010",
12234 => "11110101111101111111111011111011",
12235 => "11110110111010001110111011101010",
12236 => "11111110111101100000001011110111",
12237 => "11011010111100001111100111101101",
12238 => "00000001111101001111011000000011",
12239 => "11101001111100111111000111110010",
12240 => "11001111111100011110000011111010",
12241 => "11101101111100001101111111111110",
12242 => "11111000111011111111000111110101",
12243 => "11101111111000001110100011100110",
12244 => "11110000111101000000001111110100",
12245 => "11001011111101111110111111100100",
12246 => "11111101111010101111000111111100",
12247 => "11101100111100011110010111101010",
12248 => "11000110111011011110011111111000",
12249 => "11110100111010001100100000000010",
12250 => "11111000111010111111000111101111",
12251 => "11110001110011001110010111100000",
12252 => "11110100111011101111101011110101",
12253 => "11011011111010111111001011100100",
12254 => "11111110111010101111010011111101",
12255 => "11100000111001101101101111101110",
12256 => "10110111111011011110100011110111",
12257 => "11100101111010011100011000000010",
12258 => "11110101111010101110101111110000",
12259 => "11110000110111111111010111101100",
12260 => "11110110111100101111100111110101",
12261 => "11110101111100011111011011110110",
12262 => "11111010111011111111101100000100",
12263 => "11101111111000101110101111110100",
12264 => "11011000111110111110101011111001",
12265 => "11110010111010111101100100000000",
12266 => "11111000111110001111010011110010",
12267 => "11110100111011001111010011101100",
12268 => "00000010111111110000001111111011",
12269 => "11101110111101110000001011110100",
12270 => "00000000111101001111100000000001",
12271 => "11101101111011111111010011110110",
12272 => "11100001111101001110101000000100",
12273 => "11110100111011101110101111111110",
12274 => "11110111111100101111101011111111",
12275 => "11110101111010101111011111101100",
12276 => "11111011111110010000011011111001",
12277 => "00000000111110011111101100000000",
12278 => "11111011111110011111001111111111",
12279 => "11110101111001111110111100000010",
12280 => "11100010111101011111001111111010",
12281 => "11101010111101011110011011111011",
12282 => "11111000111110001111000111111100",
12283 => "11111011111101101111101111111010",
12284 => "11111111000000010000011011111101",
12285 => "00000110000000101111111000000000",
12286 => "11111100111110110000000011111111",
12287 => "11111111111110010000000100000101",
12288 => "11110000000000110000001011111110",
12289 => "11111100111111000000001111111011",
12290 => "11111101111111001111100100000010",
12291 => "11111101000000011111110111111110",
12292 => "00000010000000110000010000000011",
12293 => "00001101000001110000000100000001",
12294 => "11111100000001000000000100000001",
12295 => "00000011000000111111111100000110",
12296 => "11111010000000110000010000000010",
12297 => "00000010111111100000100111111110",
12298 => "11111101000001000000000100000000",
12299 => "11111101000000001111110011111110",
12300 => "00000101111111110000001000000010",
12301 => "00001000000000111111111000000000",
12302 => "00000010000000000000001111111111",
12303 => "00000000111111110000001100000110",
12304 => "11111101000000010000001111111100",
12305 => "11111111111111000001000111111111",
12306 => "00000000111111101111110011111110",
12307 => "11111001111110111111110111111011",
12308 => "11111100111111110000001011111101",
12309 => "11110101111111010000000011111001",
12310 => "11111110111110101111101100000010",
12311 => "00000011111111110000000100000001",
12312 => "11111100111111001111011100000011",
12313 => "11111110111101110000100011111100",
12314 => "11111001111110001111111000000000",
12315 => "11110001111101111111011111100101",
12316 => "11111011111011000000000011111010",
12317 => "11101011111101001111010011101101",
12318 => "00000000111010101111001011111100",
12319 => "11110000111101111111011011111101",
12320 => "11011111111000111101100011110111",
12321 => "11110101111001011110101111111101",
12322 => "11110111111010111111010111111001",
12323 => "11110011110100001111100011110011",
12324 => "11111101110110110000000111101111",
12325 => "11110111111101101111011111110110",
12326 => "11111101111011011110110111111101",
12327 => "11011010111001111111111011111011",
12328 => "11110001110111001110110111110111",
12329 => "11100101111011111110011011111101",
12330 => "11110000111011111110100011110010",
12331 => "00000011110100100000100000000101",
12332 => "11101011111100100000010111111000",
12333 => "00001011111110101110010100000100",
12334 => "11111010000001010000000011111111",
12335 => "11110001110010110000010100001101",
12336 => "00000100111110001111110011011101",
12337 => "11100101000000111111100111111111",
12338 => "11111111000010001110101111100010",
12339 => "11111100111011011111100100001001",
12340 => "11011101111100110000001000000010",
12341 => "00000010111111111110010000000011",
12342 => "11111101111101001111110111111101",
12343 => "11111100101111100000101000000000",
12344 => "00010001111111100000100111001001",
12345 => "11111100111111110001000011111011",
12346 => "00000100000000110000010111011010",
12347 => "11100100111011011111011011111101",
12348 => "11111110111101010000010100000110",
12349 => "11101001000001011110011011101101",
12350 => "00000011111101111111110011111000",
12351 => "11111111110111101111111011110110",
12352 => "00000001111100111111110011010100",
12353 => "11111000000000001111111011111011",
12354 => "00000111111101111111101011101000",
12355 => "11101110111000001111111011111001",
12356 => "11011110111100111111110111111100",
12357 => "11110000000000001110011011101000",
12358 => "11111011111110111111011011111110",
12359 => "11101110110101101111100011110000",
12360 => "11111010111100101111100011100011",
12361 => "11110010111100001111001011111010",
12362 => "00000100111101111111001011100010",
12363 => "11110000111011110000101011111111",
12364 => "11100111111110101111111011110110",
12365 => "11110010000000001111001011110101",
12366 => "11111001111101001111101100001000",
12367 => "11111000111011101111100000000100",
12368 => "11110111111010111111100011110101",
12369 => "11111100111111101111101011111111",
12370 => "00000010000000111111100111110010",
12371 => "11100101111111100000100100000010",
12372 => "11101001111100110000001011110010",
12373 => "11100100111111100000001011110000",
12374 => "00000011111110101111011000000011",
12375 => "11110101111100000000000100001011",
12376 => "00000001111011011110110011111010",
12377 => "11111111000000001111111000000001",
12378 => "00000010000000011111110111110011",
12379 => "11110010000001101111000111111110",
12380 => "11100111111010100000001111110000",
12381 => "11001011111011001111010011011110",
12382 => "00000000111001011111011000000000",
12383 => "11110000000000000000100111110101",
12384 => "00000101111101101110110111111000",
12385 => "11111011111100110000011000000000",
12386 => "11110011111100101111111111101011",
12387 => "11110011110000001111001011101100",
12388 => "11110000111111010000001011110110",
12389 => "11110001111100011111100111110111",
12390 => "11111001111100011111010111111110",
12391 => "11101010110001101101110111111001",
12392 => "10101110111101011111011011111101",
12393 => "11101011111101101100100100000010",
12394 => "11110011111101111111001011111100",
12395 => "11111011111001101111100011110011",
12396 => "00000011000000110000010011110110",
12397 => "00000100111111110000000000000011",
12398 => "11111101111111011111110000000011",
12399 => "11111100110111011111110111111111",
12400 => "11011111111110001111100111111101",
12401 => "11110011111110101110111111111101",
12402 => "11110111111101111111001000000010",
12403 => "11110000111010111111011111110111",
12404 => "11111110111100110000010011111001",
12405 => "11100111111101000000010011110100",
12406 => "00000010111101011111100100000000",
12407 => "11111010111100011111000111110100",
12408 => "11100101111100111111000000000000",
12409 => "11110110111110101111001111111011",
12410 => "11110110111110001111101100000001",
12411 => "11011110111101011110011011011011",
12412 => "11110110110110010000011011101110",
12413 => "11011000111011101111100111011110",
12414 => "11111110110111101110100100000000",
12415 => "11100000111101011110110111101110",
12416 => "11100111110101001110000011101110",
12417 => "11110001110111001101101011111101",
12418 => "11101101111001001110101011110000",
12419 => "11011101110010111110110000000110",
12420 => "11101001111101011111110111110110",
12421 => "00000011111101111101010100001001",
12422 => "11111001111001101111011111101111",
12423 => "11101110110111101111101000001000",
12424 => "11101010111110000000010010111111",
12425 => "11011010000010111111110111111010",
12426 => "11111101000001111110010011011100",
12427 => "11110001101010100000011100000100",
12428 => "11000000111110001111100000000111",
12429 => "00000000000000011100001111111100",
12430 => "11111000111001101111110011010010",
12431 => "11111101101001111111111100001001",
12432 => "11110110000000001111101010101000",
12433 => "11111010000000100000001111111100",
12434 => "00000111000000110000011011000100",
12435 => "11111011101100100000011000000101",
12436 => "00001110111101000001010000000011",
12437 => "11111111000000011111101011111111",
12438 => "11101010000001001111100011010011",
12439 => "11101111101110011111101000001000",
12440 => "11101101111110101110100011101011",
12441 => "11110000000000110000101011110101",
12442 => "00000010000001000000010111111011",
12443 => "00000010110011111111101100001011",
12444 => "00011001111110010010011100000111",
12445 => "11110110000001000001101011111011",
12446 => "11100110000010101111110111010000",
12447 => "11110001110111001111110100010101",
12448 => "11110001111110011111111011110010",
12449 => "11110101000001110000101011110100",
12450 => "11111100000010001111110100001011",
12451 => "00000110111001001111110100001001",
12452 => "00010011000000100001000000000111",
12453 => "11111010000001100001111011111100",
12454 => "11110101000011000000000111110011",
12455 => "11111111111000010000101100001101",
12456 => "11111110000001010000100100010001",
12457 => "11110000000100000000110011101010",
12458 => "00001001000010001111011100001010",
12459 => "11111011111011000000101000001100",
12460 => "00010010000000110000010100001011",
12461 => "11111010000011110001100011110001",
12462 => "11110110000001010000000100001001",
12463 => "11111011110001110000111000010001",
12464 => "00000011000001000000000100010010",
12465 => "11111001000001110001011111100100",
12466 => "00001111000000011111110000010000",
12467 => "00000010000001110000011000000100",
12468 => "00010010000001110001100000000111",
12469 => "11100011000101110001111011011101",
12470 => "00000010000010000000000000010001",
12471 => "11111000111100000000110100000101",
12472 => "00010010111101111111110000010101",
12473 => "11110111111110010000110011111001",
12474 => "00001110111101110000011100011100",
12475 => "00001101000001011111110111111110",
12476 => "11111000000011011110100011110111",
12477 => "11101110000001000000000011100000",
12478 => "00000110000100000000101111110001",
12479 => "11111011111001100000011111101111",
12480 => "00000111111010110000000100001100",
12481 => "11111110111111110000101011111011",
12482 => "00000110111101011111101100000110",
12483 => "11111000000000010000110111110001",
12484 => "11001100000000111101000111110111",
12485 => "11101011111111001010110011101110",
12486 => "00000010000000000000001100000001",
12487 => "11111111111111100000010111110101",
12488 => "00001100111101000000010011001110",
12489 => "11111110111110101111111111111010",
12490 => "00000000111111011111011111001110",
12491 => "11110001111101111111111000000001",
12492 => "10111011111000111110000111111000",
12493 => "11011100111101111011111011101001",
12494 => "11111111111100101111100100000101",
12495 => "11101010110111011111011100000100",
12496 => "11110111111001101110011011101100",
12497 => "11110010111100001111101100000010",
12498 => "00000000111100000000000111011010",
12499 => "11110001111101101111000011110101",
12500 => "11011100111101101111101011110101",
12501 => "11100111110111101110101111110000",
12502 => "11111100111001011110111011111101",
12503 => "11100110111010100000011011101100",
12504 => "11110010111100101110111011111011",
12505 => "11101101111010100000000011111011",
12506 => "11110100111011001111000111101111",
12507 => "11110011111000001111000011101000",
12508 => "11011111111011101111110111110001",
12509 => "11101111111011111110001111101111",
12510 => "11111010111101101110111111110101",
12511 => "11110110110111001110111011111010",
12512 => "11010010111000001111011011100111",
12513 => "11101111111010111110001000000001",
12514 => "11101110111100011111000011101001",
12515 => "11011001111000101111000011110011",
12516 => "11000110111001110000000011110100",
12517 => "00001000111100001011111011111110",
12518 => "11111101110110101111001011100011",
12519 => "11100100111000111111110000001010",
12520 => "11010101111011111111000011001000",
12521 => "11101111111110101111000111111111",
12522 => "11110110111100111111001011001110",
12523 => "11101111110011110000001000000010",
12524 => "11101011111001100000100000000110",
12525 => "00000001111111011110001100000011",
12526 => "11110111111100101111010111101010",
12527 => "00000011111101011111100100000011",
12528 => "11011100111110111111110111100001",
12529 => "11111001111101110000101011111001",
12530 => "11111001111111100000000011011100",
12531 => "11110011111001111111110000000111",
12532 => "00010100111000110001110000000001",
12533 => "00000100000000001111101100000111",
12534 => "11011001111100111111011011011010",
12535 => "00001100000110001111000000011000",
12536 => "11010110111111001111101011110001",
12537 => "00001101000000010000010011111000",
12538 => "11111011111111110000101011101110",
12539 => "11111110111011011111011100010010",
12540 => "00011011111100010011010000000101",
12541 => "11111110111111110001010100000001",
12542 => "10101110111111101111100011001010",
12543 => "11110110001000111111001100100000",
12544 => "11001110111111101111101011111001",
12545 => "11111011000000000001011111101111",
12546 => "00000010000001010000010011111100",
12547 => "11111111111100011111010000001110",
12548 => "00010001111101110001101100000110",
12549 => "00000110000000100001011100001101",
12550 => "10100111000000001111110111001111",
12551 => "11111001000100100000010100101100",
12552 => "11100000111111111111101111111101",
12553 => "11111101000000110001101111011100",
12554 => "00000011000000110000001111111110",
12555 => "00010110111101100000010100001101",
12556 => "00001010001000000000010000000111",
12557 => "11111101000011010010000000001001",
12558 => "11101110000110110000101111111001",
12559 => "00001100000000010001001000100011",
12560 => "11111000000001110001111000011001",
12561 => "00001001000011100010111011000111",
12562 => "00001010000100000000100000001011",
12563 => "00001000000001110000101011111101",
12564 => "00001110000101110000001100001001",
12565 => "00000010000001110001110111110011",
12566 => "00010001000011000000100011111011",
12567 => "00001100111110110001011000001000",
12568 => "00011000000000010000111100001110",
12569 => "00000101000011010001100011010001",
12570 => "00000010000010010000000000010000",
12571 => "00001100000010010000100111110101",
12572 => "00000110000011111111110111111110",
12573 => "11111100111110100001010111101011",
12574 => "00001101000010100000010100000111",
12575 => "00001001111111110000100111101110",
12576 => "00010001111111100001001100001101",
12577 => "00000011000011000000101111101000",
12578 => "00000000000010101111100100001000",
12579 => "00000000000001110000010111111001",
12580 => "11111011111111111110000011111100",
12581 => "11110010111101000000100111100111",
12582 => "00001001111111100000000000001101",
12583 => "11111111111100000000101111100101",
12584 => "00010000111111011111101100010000",
12585 => "11111111111111001111111111110100",
12586 => "11111100111111101111111100000001",
12587 => "11111100000000101111011111110110",
12588 => "11111110000000111110101111111001",
12589 => "11011101000000000000010111011111",
12590 => "00001001000001011111110100011110",
12591 => "11111111111101000000100011000000",
12592 => "00000111111101000000001100010101",
12593 => "11111010111110001111110011110111",
12594 => "11111110111101110000011000001010",
12595 => "00000000111110101111110011110110",
12596 => "11110000000010001110110111110011",
12597 => "11001001000000001110010011011101",
12598 => "00000100111111010000101100010001",
12599 => "11101111111101100000000011001010",
12600 => "11111100111010111111110111110011",
12601 => "11110101111111001111011000000000",
12602 => "00000101111101011111010011110100",
12603 => "11111010111111111111001011100010",
12604 => "11110100000000001111100011101100",
12605 => "11101111111100101110111111111000",
12606 => "00000000111101011110110100000010",
12607 => "11101100000000001111110111011010",
12608 => "11111100111100000000000111111011",
12609 => "11110000111100011111100000000000",
12610 => "11110101111100101111000111101101",
12611 => "11111110111001101111001111111000",
12612 => "11010000000000111111100011111100",
12613 => "11111110111100101101100011111101",
12614 => "00000000111110001111100011111010",
12615 => "11110000111000111111100000000100",
12616 => "11101100111110001111110011110111",
12617 => "11110010111111011110101000000010",
12618 => "11111000111110011111000111010101",
12619 => "11110011000100011111011100001100",
12620 => "11011101111101111111101000000111",
12621 => "00010011000001011101110000001100",
12622 => "11111111111110001111100111110111",
12623 => "11111101000011101111011000001010",
12624 => "11110111000001110000001011111011",
12625 => "00000001000001000000011100000001",
12626 => "11111001000010100000000011011011",
12627 => "00000001000001001111110100001001",
12628 => "00000111111111000001001100000010",
12629 => "00000100111111111111101000000111",
12630 => "11101011000010010000010111101100",
12631 => "00000101000101101111101100010011",
12632 => "11011010000000010000100111111000",
12633 => "11111101000001000000110011110111",
12634 => "00000100000000100000000011110111",
12635 => "00001011000100110000100000001011",
12636 => "11111110000001110000010100000101",
12637 => "00000110111111100000000000001011",
12638 => "11011000000010100000010111011100",
12639 => "00001110000101111110110100001000",
12640 => "11011101000010110000111111111110",
12641 => "00000111000011000000111111101110",
12642 => "11111111000001100000010011110111",
12643 => "00001010000010010000111100000110",
12644 => "00000001000010001111100100000101",
12645 => "00010011000010001111100000001101",
12646 => "11000001000010010000011111011100",
12647 => "00000111000100011110111000011010",
12648 => "11101100000010100000110100000011",
12649 => "00000001000001000000001111100110",
12650 => "00000111000010010000000100000010",
12651 => "00001100000001110000101011111111",
12652 => "00001110000101111111111111111110",
12653 => "00010100111111000000000100010100",
12654 => "11001100000100000000000111110101",
12655 => "00010000000001100000010000101100",
12656 => "11111010000010110001001000000110",
12657 => "00010001000101010000111011001001",
12658 => "11111111000100010000110011111111",
12659 => "00001111000000110001010011111111",
12660 => "00000110000101010000001100010000",
12661 => "00001010000011010000011100010111",
12662 => "11010100000100100000001111111100",
12663 => "00010110000001100000101000100000",
12664 => "00000011000010010001101100000101",
12665 => "00010111000100010001101010110011",
12666 => "11111101000101010000111000000000",
12667 => "00000011000010100000110111111100",
12668 => "00000000000100110000010000001100",
12669 => "11101100000001000000011011110001",
12670 => "11111110000010000000011011100110",
12671 => "00001011000010011111101000010111",
12672 => "00000101111101110001001011111001",
12673 => "00001011000011100001001111001001",
12674 => "00000110000010100000001100000011",
12675 => "00000000000010000000101111111011",
12676 => "00000001000000101111101100001011",
12677 => "11111000111111000000000111111110",
12678 => "00001111000000010000001111111110",
12679 => "11111100111111100000000000001001",
12680 => "00000100000001010000011111110111",
12681 => "11110110000010010001001111100100",
12682 => "00000001000001100000100100000011",
12683 => "11111001000000100000001111101100",
12684 => "00000011000001001111010100000000",
12685 => "11100110111101100000001011100110",
12686 => "11111010000001110000001111111110",
12687 => "11111011111101011111110111101011",
12688 => "00010001111101000000000111111110",
12689 => "11111110000010100000000011101101",
12690 => "00000111111101100000000100000101",
12691 => "00000001000010100000000111110110",
12692 => "11111100000001111110101111110111",
12693 => "11011100111111001111010111101011",
12694 => "00000100111111100000000100001011",
12695 => "00000101111110100000111011101101",
12696 => "00010010111010100000100111111001",
12697 => "11111100000010100000100000000111",
12698 => "00000000111110110000000100000001",
12699 => "11111010000000011111001011111010",
12700 => "11101101111101101110111111110011",
12701 => "11111010111011101110011100001000",
12702 => "00000100111100101111110000001001",
12703 => "11111010111101110000110011101101",
12704 => "00001001111101111111010111110011",
12705 => "11111011111011010000001100000011",
12706 => "11110010111101101111011011101100",
12707 => "11101010111110011111010111111000",
12708 => "11100100111001101110111111110011",
12709 => "00000100111000001110011111111101",
12710 => "11111111110111111111010011111010",
12711 => "11110100111100101110100100000000",
12712 => "11101111111100111110001111100101",
12713 => "11111111111011101110101000000000",
12714 => "11110001111011111111110011100000",
12715 => "11110011111100001111100111111111",
12716 => "11111111000000011111111111111011",
12717 => "00001000111101101111101000000101",
12718 => "11111110111111001111111011111110",
12719 => "11110100111101111111010011111110",
12720 => "11110011000000101110110100000101",
12721 => "11110001111110011110111011111110",
12722 => "11110111000000101111001111111011",
12723 => "00000110001010000000011000001010",
12724 => "11110011000010111110000000001001",
12725 => "00001101000010101111001000010011",
12726 => "11111000000001010000001011111100",
12727 => "00001010000111111111111100000000",
12728 => "00000110000010000001011011111010",
12729 => "00001101000010100000101011111111",
12730 => "00000110000001110000100011110011",
12731 => "00001101000110110000010100001010",
12732 => "00001001000011011111111100000101",
12733 => "00001100000001010000101100001011",
12734 => "11110001000011000000010111110011",
12735 => "11111101001000101111101000000011",
12736 => "11111001000000110000111111111111",
12737 => "11111110000011000000100011110100",
12738 => "00000011000010010000001100001000",
12739 => "00001111000111100000110111111111",
12740 => "11111001000101101110010100001100",
12741 => "00001000000000111111010100000101",
12742 => "11110001000010000000101011101100",
12743 => "00010011000011011110000111100111",
12744 => "00001111000001100001011011111100",
12745 => "00001000000010100000010011100111",
12746 => "00001010000001100000011011111111",
12747 => "00010000000100110000001111110100",
12748 => "00000111001000001110100000000111",
12749 => "00001010000010011111110000000110",
12750 => "11110100000100110000101000001001",
12751 => "11111111111110101111100111101010",
12752 => "00010011000010110001001100010011",
12753 => "00000111000011010000010011001101",
12754 => "00001011111111110000011000000010",
12755 => "00001111000010000000110011110010",
12756 => "00000111000111111111011100000001",
12757 => "11111100000011100000010100000101",
12758 => "11101001000010111111111000011110",
12759 => "00001110000001001111110111110110",
12760 => "00010111000000100001010100011010",
12761 => "00001100000001010000111011000110",
12762 => "00000110000010000000111000001101",
12763 => "00010111111010110000100100001010",
12764 => "00010111000100000000101100001001",
12765 => "11110101000100100001000111111111",
12766 => "11001101000101100000011000001000",
12767 => "11111100000010001111110100011100",
12768 => "11111011111111100000110000010100",
12769 => "11111111000101010001001111011001",
12770 => "00000111000101000000001000001110",
12771 => "00001101111000100000111100001110",
12772 => "11110101111111101101100100001001",
12773 => "11100101000010011111101111110001",
12774 => "11011100000010010001010111101000",
12775 => "00000101111010100001000000001111",
12776 => "11110100111110010001000011110111",
12777 => "00001001000101100001111111100111",
12778 => "00001001000010000000100111111100",
12779 => "11111111000001011111111111111111",
12780 => "00000111000000011111001000000101",
12781 => "11101001111111110000100111110011",
12782 => "00000110000010000000101000000000",
12783 => "11111011111111100000000111110011",
12784 => "00001000111111101111111011111000",
12785 => "11110110000000001111111011101000",
12786 => "00001101111111010000010000010010",
12787 => "11111001000001100000001011110111",
12788 => "11101110111111111110000011111101",
12789 => "11101100111111001110011011101100",
12790 => "00000000000000000000110000000000",
12791 => "11111011111110101111010011101010",
12792 => "00010001111100011111101011110011",
12793 => "11111010000000001111001111110000",
12794 => "00001000111101111111111111111111",
12795 => "00000011111111110000000011110111",
12796 => "11110000000010011110011011111001",
12797 => "11101111111111011110000111110111",
12798 => "11111000111111110000101011111001",
12799 => "00010001111111111110000111010111",
12800 => "00001001111101010000101011110010",
12801 => "00000111000001001101111111110111",
12802 => "00000110000000010000000011101101",
12803 => "00000011000010101111111111110010",
12804 => "11111110000000101111110011110111",
12805 => "00000010111111001111011000001010",
12806 => "00000001000000000000010100001000",
12807 => "00000010000001001111001111100010",
12808 => "00010100111110110000100111111101",
12809 => "00000001111111001110001111111111",
12810 => "00001000111011110000000000000100",
12811 => "11111001111110111110110011100010",
12812 => "11101100000000111111100011110000",
12813 => "11111101111010111111001100000010",
12814 => "11111011000010011111000111110111",
12815 => "11110111111110111111100011101111",
12816 => "11110001111110111111101011110010",
12817 => "11111000111110011110100100000001",
12818 => "11111000111010111111001011110001",
12819 => "00000001111110111111100111111111",
12820 => "11110010111111101111101111111011",
12821 => "00000010111110011111101000000010",
12822 => "11111111000000011111111111111111",
12823 => "11110111111100101111000111110110",
12824 => "11110101000000011111001000000011",
12825 => "11110001000000011110111100000000",
12826 => "11111111000001101111101111110011",
12827 => "00001101000111010001001100000110",
12828 => "11111101000101001110110000000110",
12829 => "11111111000011000000010000000101",
12830 => "11111010000000110000000100000000",
12831 => "00001111000100101110100011101001",
12832 => "00001011000001000001011000000000",
12833 => "00010010000001110000001111110010",
12834 => "00000000000000110001000000000011",
12835 => "00001010001000010000001000000011",
12836 => "00000011000100011111011100000001",
12837 => "00000010111110100000001000000000",
12838 => "00000010000011100000011000000011",
12839 => "00000001000010101110000011101101",
12840 => "00000100000000110000000100000110",
12841 => "00000001000001111111111111111010",
12842 => "00000100000001010000011000000100",
12843 => "00001010000111110000001111111001",
12844 => "11110111000101111101110100000111",
12845 => "11111111000000101111011000000000",
12846 => "00000001000000110000000011111110",
12847 => "00001000111101001110111011010000",
12848 => "00010011111111100000111100000001",
12849 => "00001110000000111111011011110010",
12850 => "00000100000000010000100100000010",
12851 => "00000000000010100000001111111011",
12852 => "11101111000011111110001011111011",
12853 => "11111101111110011111110011110100",
12854 => "00001011111110111111110100011101",
12855 => "00000011111101100000000011001111",
12856 => "00011010000001010000100000001010",
12857 => "00000010111111101111100111010101",
12858 => "00000000111111110000101011111011",
12859 => "00000001111100010000100111111100",
12860 => "11111100000010011111010011111000",
12861 => "11101000000000110000111111101000",
12862 => "11110001000000001111111000101100",
12863 => "00001010111100001111101011101100",
12864 => "00001111000000100000011100001101",
12865 => "00000111111110100000010011010101",
12866 => "00000011000000110000000100001001",
12867 => "00010100101111100000011100000111",
12868 => "00011010000001010001001100001101",
12869 => "11110010000010100001111011111100",
12870 => "11001101000100110000100100001000",
12871 => "00000100111101010000011000100010",
12872 => "11111000111111110000111100011101",
12873 => "00000110000010110001101111100100",
12874 => "00001000000011100000001100000110",
12875 => "00010011111011100000111100000011",
12876 => "11111001000001011110100111111111",
12877 => "11011111000001100000011011100100",
12878 => "11010101000100100001001100000001",
12879 => "00010010000001100000010000000001",
12880 => "11101101111101010000110000010011",
12881 => "00001000000000101111111011010111",
12882 => "00001101111111110000000100001011",
12883 => "11111101000001010000000100000110",
12884 => "11101101111010001110011000000110",
12885 => "11101100000000011101000111101010",
12886 => "11011011111111010000111011100000",
12887 => "11111110000001011101111011101100",
12888 => "11101111111101001111100011100001",
12889 => "11111101111111101110000111111110",
12890 => "00001010111111001111110111100000",
12891 => "00000110000001000000010000000001",
12892 => "11110100111110101111000100000100",
12893 => "11111010111110011110101100000011",
12894 => "11110011111110000000101011011010",
12895 => "00001001000001101110001111111111",
12896 => "11100111111111011111011111110011",
12897 => "00000110000001011110011011110101",
12898 => "00000001000000010000101011101111",
12899 => "00000001000011101111111100000000",
12900 => "11111101111100111111110011111111",
12901 => "11111010111111001110011000000011",
12902 => "11110110111110010000010011011000",
12903 => "00000100000011011101011111110100",
12904 => "11101101111101111111111011100011",
12905 => "00000010111111001101101011111001",
12906 => "11111111000000011111110111110111",
12907 => "00000100000000011111010011110000",
12908 => "11111101111100011111110011101111",
12909 => "11100001110110101111011111101111",
12910 => "11110011111101100000001111110110",
12911 => "11111101000001011100111011111000",
12912 => "11101001111011101111111011111110",
12913 => "11111010000000001100011011111101",
12914 => "00000010111001111111111000000100",
12915 => "11100110111000111110100011101101",
12916 => "11101010111011101111110011101011",
12917 => "00001001111001101110011111111110",
12918 => "11111101111001101110110111111011",
12919 => "11101110111001011110101000000110",
12920 => "11011111111101001101101111100011",
12921 => "11101000111000001100001111111111",
12922 => "11110000111011101110101111011110",
12923 => "00000001111111000000000100000010",
12924 => "11101101111110100000001011111111",
12925 => "11110111000000001111000111111100",
12926 => "00000000000001001111111011110111",
12927 => "11111000111110001111101011101101",
12928 => "11101101111111101110101111111100",
12929 => "11111001111111101111010000000000",
12930 => "11111101000010000000000011101011",
12931 => "00001110000010110000010111111010",
12932 => "11111110000010011111101111111111",
12933 => "11111010000000010000001011111000",
12934 => "11111110111110110000000111111100",
12935 => "00000101111110101101100011100110",
12936 => "11111010111110110000111000000110",
12937 => "00000001111111111101100011111001",
12938 => "00000001000001000000001000000111",
12939 => "11111110001000001111100100000101",
12940 => "00000101000010101110111100000101",
12941 => "11110111000000000000000011110111",
12942 => "00000011000001111111101000000011",
12943 => "11110101111101101110101111010111",
12944 => "00010111111111010000000000001100",
12945 => "00001000111111000000011011111000",
12946 => "00000000000001010000010000000111",
12947 => "11111100000011101111100111111101",
12948 => "11111010000001001101101011111110",
12949 => "11101100000001001111011011110100",
12950 => "00001101111111101111101000001000",
12951 => "11110001111010011110101011001111",
12952 => "00011001111110000000001000001001",
12953 => "00000111111101101110110011110001",
12954 => "11111101000000101111111000000000",
12955 => "11111011111101110000011000000010",
12956 => "11111111000011001110011111111010",
12957 => "11101000000001110000010011100100",
12958 => "00001100000000111111101100100101",
12959 => "00000011111000100010001011011111",
12960 => "00101011000000010000010100010000",
12961 => "00000111111101000000100011011101",
12962 => "11111101111110010000000100001110",
12963 => "00001111110111100000011000000001",
12964 => "00011000000010100001001111111101",
12965 => "11011001000100100010010011010000",
12966 => "11110110000011100000010000100000",
12967 => "00000101111100110001111100011110",
12968 => "00011110111011100000100000010110",
12969 => "11111111000010000001101011010100",
12970 => "00000011000000000000001100010111",
12971 => "00010000101111010000101111111011",
12972 => "00010100000000100001011000000000",
12973 => "11101101000001010001101011111110",
12974 => "11100100000101100000001111110110",
12975 => "00000110000001010000110100100100",
12976 => "11110011111100010000101100001101",
12977 => "11101111000010000001001011101110",
12978 => "11111110000010010000010000000001",
12979 => "00000000111100110000110111111101",
12980 => "00000010111100110000010111111100",
12981 => "11110110111111010000101111111000",
12982 => "11011101000000100000101000000011",
12983 => "00001101000010111111000011111001",
12984 => "11100010111110110000110000001010",
12985 => "00001010000010111110011111100111",
12986 => "11111011000001000000010000001001",
12987 => "00001001000011000000011100000110",
12988 => "11111011000000011111111000000001",
12989 => "11111010111101011110110000000001",
12990 => "11001101000000100000011011011001",
12991 => "00000101000010111100011000010000",
12992 => "11100011111110110000100011110001",
12993 => "11111001000011101101111011111010",
12994 => "00000001111111100000101111110111",
12995 => "00000110000001110000010000000011",
12996 => "11111010111100111111101111111110",
12997 => "11111101111101001110101000001000",
12998 => "11101010111110000000000011100011",
12999 => "00000001000011001101110111111010",
13000 => "11011101111110111111110111110000",
13001 => "00001000000001011110011111111010",
13002 => "00000000000010100000011111110010",
13003 => "11111110000100011111101011110001",
13004 => "11111111111110100000001011111010",
13005 => "11111100111011011110111000001001",
13006 => "11111010111111011111110111110110",
13007 => "00000000000100101101111000000000",
13008 => "11110001111101101111010111110010",
13009 => "11110111111110001101111000000011",
13010 => "00000001000000011111110111111011",
13011 => "11101111000000001110101011101100",
13012 => "11101011111000001111011011101100",
13013 => "11100100111010111101111011111110",
13014 => "11111100111011011110101111111100",
13015 => "11110010000000111110100011111010",
13016 => "11110101111001101110000111101101",
13017 => "11110101111000111101111100000001",
13018 => "11110101111100001111010111100111",
13019 => "11101010110011101110101111101100",
13020 => "11010111111100011110111111101010",
13021 => "11111011110111101101111111111101",
13022 => "11111110110111001110101000000100",
13023 => "11101010110010011110000011111000",
13024 => "11001111111101011110011111101001",
13025 => "11101010111010011100110011111011",
13026 => "11101001111101001110101111011101",
13027 => "00000000111011101111110111111000",
13028 => "11101011111100000000000011111100",
13029 => "11110101111111001110101111111001",
13030 => "11111110111111011111111011111101",
13031 => "11111101111011111111001011101110",
13032 => "11101000111111111111000011111101",
13033 => "11111101111100111110100111111111",
13034 => "11111010000000001111110011101101",
13035 => "11110011111000111111011111110111",
13036 => "11110010111110011111110000000001",
13037 => "11111000111110111111101111110111",
13038 => "00000100111111001111111011111111",
13039 => "11110111110101101101100011101101",
13040 => "11001010111111101111001111110110",
13041 => "11110110111100011101101000000100",
13042 => "11111111111111100000000011110101",
13043 => "00000001000010000000000011110011",
13044 => "11111101111101111111010011111100",
13045 => "11110010111101111111101011110010",
13046 => "00001000111110001111111000000011",
13047 => "11111001111010101111000111100110",
13048 => "00001000111101001111111000000111",
13049 => "11111100111111101110101111111010",
13050 => "11111010111110101111010100000100",
13051 => "11111011111101110000001111101100",
13052 => "00000011000000111111011011111010",
13053 => "11011110111111100000001111100010",
13054 => "00010000000000111111101000000110",
13055 => "11110001110110111111111011001101",
13056 => "00010010111110111111110000001001",
13057 => "11110010111101001111001011111001",
13058 => "11111110111101101111101100001100",
13059 => "11111101111000110000011011110111",
13060 => "00010100000101101111111111110000",
13061 => "11010110000001100001011111010101",
13062 => "00001110000000101111101100011101",
13063 => "11111010110000010001111111110111",
13064 => "00101111111110100000010000010011",
13065 => "11111001000000100000001111101111",
13066 => "00000101111110001111100100011011",
13067 => "00000101110011100000000011111111",
13068 => "00001101000000000001011000000000",
13069 => "11011110000001010001110011100100",
13070 => "11111111000001001111111100000011",
13071 => "11101000111010010010001100010001",
13072 => "00010001111100011111010100001010",
13073 => "11110000000000010001101011110001",
13074 => "11111001111111011111101000010011",
13075 => "11111100111010011111101111110100",
13076 => "00001101000000010000101011111011",
13077 => "11110110000000111111111100000010",
13078 => "11110010000001001111111011110111",
13079 => "00000011111110101111001100001101",
13080 => "11010010111110110000001000001001",
13081 => "11111110111111011111010111111110",
13082 => "11111011000000110000000011111001",
13083 => "11111110111101010000000011111110",
13084 => "11111101111101001111110111110011",
13085 => "00000001111110011111101100001000",
13086 => "11011011111110111111111111111100",
13087 => "00000000000001111110111100001010",
13088 => "11100100111111000000001000000000",
13089 => "00000010111111111110100011101101",
13090 => "11111100111111011111011111110001",
13091 => "11111111111111000000001011111000",
13092 => "11101111111111001111000011111100",
13093 => "00000011000000111110111000000110",
13094 => "11100001111111110000011011110111",
13095 => "00000011000010011010101011111111",
13096 => "11010110111110111111111011110111",
13097 => "00000001000000011100001011111011",
13098 => "11111110000001001111101011110001",
13099 => "11110111000000100000000011101111",
13100 => "11100100111111011110101011110111",
13101 => "00000001111111111101011111111011",
13102 => "11101000111111010000000111101000",
13103 => "00001011000001011100001111110100",
13104 => "11100000000000001111111111011010",
13105 => "00000000111110101100011000000010",
13106 => "11111111000000010000001011011110",
13107 => "11110100000010000000000111110000",
13108 => "11111001111010101111011111111000",
13109 => "00000101111011101110100011111111",
13110 => "11111010111001111111011000000011",
13111 => "00000010000011001111000000000000",
13112 => "11111101000001001111100011101000",
13113 => "11111011111101111110110111111111",
13114 => "11101111111011001111110111110011",
13115 => "11101011111110011110111011111101",
13116 => "11100100111010111111001111101101",
13117 => "00000100111100001110010011110111",
13118 => "00000111111001011110110100000100",
13119 => "11110011111111001111101100001111",
13120 => "11111001111110011111000111100111",
13121 => "11111010111100011111101100000011",
13122 => "11101000111011101110111011100111",
13123 => "11101110110111111111010111110001",
13124 => "11000101111011101110000111101111",
13125 => "11111100111001001100010100000011",
13126 => "00000000111001001110111000000001",
13127 => "11110111110101111111001011101110",
13128 => "11101011111100111111000011101100",
13129 => "11111001111010111110111100000001",
13130 => "11101101111101111111010011011110",
13131 => "11111001111011101111110111101100",
13132 => "11100110111001001111100011111001",
13133 => "11101001111000011110011011110010",
13134 => "00000000111100111111010111110011",
13135 => "11111101111010111110111111100110",
13136 => "11101000111101101101111011110111",
13137 => "11110111111010111110111011111111",
13138 => "11110010111100111111010111110101",
13139 => "11110111111101011111100111110111",
13140 => "11110000111101111110110111111010",
13141 => "00000011111101011111000000000001",
13142 => "11111110111110111111110111111000",
13143 => "11111001111011001111000100000001",
13144 => "11101110000001011111101011110111",
13145 => "11110110000000001101110111111101",
13146 => "11111100000000011111101111110001",
13147 => "11110110000011011111100011110000",
13148 => "11110101111100101111011111111010",
13149 => "11101101111011111111101111110000",
13150 => "11111111111110111111101011111110",
13151 => "11111100111110101111011111101110",
13152 => "00000100111011011111000111110111",
13153 => "00000110111100111111000100000100",
13154 => "11110101111011011111101111111010",
13155 => "11111011111101001111100111110101",
13156 => "00000100111110100000100111101110",
13157 => "11110111111101000000101111110101",
13158 => "00010011111101111111010100001110",
13159 => "11101101111010100001101000001000",
13160 => "00010110111101111111100100000001",
13161 => "11101100111111100000011000000011",
13162 => "11110010111100111111010100001011",
13163 => "11111110110010101111101011111011",
13164 => "00010010111110010000101011110111",
13165 => "11101000111011110001010111110000",
13166 => "00001010111100001111101000001111",
13167 => "11110100101110110001101000001000",
13168 => "00001011111101011111001000001110",
13169 => "11101110111111100000110000000001",
13170 => "11111001111101101111100100010111",
13171 => "11110111110110101111001111110110",
13172 => "00010011111110110001101011111000",
13173 => "11101101111101110001000111101011",
13174 => "00000111111111011111010011101101",
13175 => "11100110111110100000010000010100",
13176 => "11110011111011011110100100000000",
13177 => "11100111111101111111111100001010",
13178 => "11111011111101111111011100001001",
13179 => "11110001000001011111000011111100",
13180 => "00000000111010100001010100000000",
13181 => "00001010111111001111011000001010",
13182 => "11111100111100111111011011110000",
13183 => "11111110000011110000000000010100",
13184 => "11111000000010011111011111110011",
13185 => "00001000111011011111110100000001",
13186 => "11101101111110111111110111110111",
13187 => "00000000111111011111111011111010",
13188 => "11101100111011111111110111110111",
13189 => "00000101111111111110001000001111",
13190 => "11111011111101011111111111111100",
13191 => "11111001000001111111010100000111",
13192 => "11101100000000111111110111110111",
13193 => "11110111111111011110100000010110",
13194 => "11110011000000011111000111100101",
13195 => "11111010111110101111110111111110",
13196 => "11101010111101111110011111111000",
13197 => "00000111111101001110011000000110",
13198 => "11110010111010100000000111110111",
13199 => "11111100000000001100110111111101",
13200 => "11101101111111101111110111111011",
13201 => "11111111000000011101001000000001",
13202 => "11111001111111011111111111100101",
13203 => "11111100111110010000010111111110",
13204 => "11110100111110111110100000000001",
13205 => "00000011000001101110110000001010",
13206 => "11101111000000110000000111110111",
13207 => "00001100111111001101111011111000",
13208 => "11111000000010000000101111101110",
13209 => "00000000111111011101110011110010",
13210 => "00000001000001000000000011110000",
13211 => "11110101000000011110111111111000",
13212 => "11110000111110101110111111111001",
13213 => "00001000000000111110110100000001",
13214 => "11110111111100001111111011111011",
13215 => "00000000000001011111010000000100",
13216 => "11111110000000011111110111110101",
13217 => "00000001111110001110110011111110",
13218 => "11110111111101101111010011110101",
13219 => "11111011111111010000010000000010",
13220 => "11110100000000011111001111110101",
13221 => "00010011000001101111001000001111",
13222 => "11111111111100111111111000001101",
13223 => "00000110111101100001001100001001",
13224 => "00001010000010000000010111110111",
13225 => "00000100000000100000000111111001",
13226 => "11111110000010101111001111110110",
13227 => "11110100000000001111101000001010",
13228 => "11110010000000101111001011111111",
13229 => "11111000000010101101100000000000",
13230 => "11111111111111101111110111111100",
13231 => "11111101111101010001000011101001",
13232 => "00010001000000101111100111101001",
13233 => "11111101111100100001001111111111",
13234 => "00000010111111001111011011101011",
13235 => "11110001000000101111100111111100",
13236 => "11100010111100101111100011110010",
13237 => "11110010111110101101111111110100",
13238 => "11111010111101111111010111110100",
13239 => "11110101111111010000000100001000",
13240 => "11110111111100101111000011101001",
13241 => "11111001111110101111001100000010",
13242 => "11111100111101101111010111011101",
13243 => "11110111111011111111011111110010",
13244 => "11111110111010001111111011111101",
13245 => "00000100111100100000000100000011",
13246 => "00000011111100001111110100001001",
13247 => "11110110111101101111101111110111",
13248 => "11111111000001101110110011111111",
13249 => "00000100111100101111011100000010",
13250 => "11111001111100111111111000000001",
13251 => "11110111111101011111000011110111",
13252 => "00000001000011001111110111110100",
13253 => "11110010111111010000000011110100",
13254 => "00000010111111101111101111111110",
13255 => "11110100111010101111101111111110",
13256 => "00001011111101011111110111111100",
13257 => "11110111111111001111000000000100",
13258 => "11111110111101011111001000000000",
13259 => "11101111110011111110111000000111",
13260 => "00000000111111110000110111111111",
13261 => "00000000000010011111111111111110",
13262 => "00000010111111001111100111111110",
13263 => "11110000110101000001100000011011",
13264 => "11111101111111111110111111110011",
13265 => "11101110111110100000110111111101",
13266 => "00000001111110000000000000000010",
13267 => "11110001111100011110111000000000",
13268 => "00010011111101110001110011111101",
13269 => "11110111000000000000110011111000",
13270 => "00000100111110011111001111101000",
13271 => "11111000111010010001101000001011",
13272 => "00001000111101011110111111111010",
13273 => "11110110111011000000101000000101",
13274 => "11111001111100101111111000010001",
13275 => "11110010111111001111010000001001",
13276 => "00000100111101100000111000000001",
13277 => "00000010111101001111100100000111",
13278 => "11111001111101001111100111011101",
13279 => "11101110111111010001001000010111",
13280 => "00000101000000101110110011110001",
13281 => "11111000111110010000101100001100",
13282 => "11110111111111001111110111111110",
13283 => "11101111000010101110110111111010",
13284 => "11101110111100101111100111111000",
13285 => "00000011000000101101100000000011",
13286 => "11111101111100001111001111110101",
13287 => "11111001000000100000011000001001",
13288 => "00001010000000111111011011101100",
13289 => "00000000111010101111100011111110",
13290 => "11110110111101011111011111100111",
13291 => "11101000111111111111101000000001",
13292 => "11110100111010011110111011111100",
13293 => "00001001111111001101011100000101",
13294 => "11111110111011101111010011110110",
13295 => "00000101111111010000001011111101",
13296 => "11111111000000101111100011101011",
13297 => "00000001111010101111001000000010",
13298 => "11111000111111000000001111100101",
13299 => "11110001000000101111110100000010",
13300 => "11111010111011011111110011111100",
13301 => "11111110111111011111000011111111",
13302 => "11101101111110001111111111110111",
13303 => "11111000000000101110100111110011",
13304 => "11111100000000011110100111110101",
13305 => "11111011111011011110110100000101",
13306 => "11111010111110011111101111111001",
13307 => "00000000111111111111100111111101",
13308 => "11111100111101111111100000000001",
13309 => "00001010111110111111110000001001",
13310 => "11110010111101011111110000001011",
13311 => "11111010000000101110110011101100",
13312 => "11111100000010110000010100001011",
13313 => "11111010000000101110110100000000",
13314 => "11111011000000011111100000000000",
13315 => "00000011000011001111111111110010",
13316 => "11110111000001001110010111110101",
13317 => "11111110111100011111001100000000",
13318 => "00000011000000111111110000001111",
13319 => "11111001111111010000011011011110",
13320 => "00001111111111011111011111111100",
13321 => "00000000111111010000001011111011",
13322 => "00000000000000001111111011111000",
13323 => "00000000000001110000010000000000",
13324 => "00001010000001110000010100000100",
13325 => "00010011111111110000111000010100",
13326 => "00000011000000100000011000010101",
13327 => "00000110111111000000111100000000",
13328 => "00001110000100000001000100010001",
13329 => "00000001000000110001100000000000",
13330 => "11111101000010000000010100001010",
13331 => "00001000000011000000101000000010",
13332 => "00001010000000000000011000000101",
13333 => "11111010111110000000101111111010",
13334 => "00000011000000110000001100000011",
13335 => "11111011000011011111111011111101",
13336 => "00001000111110110000101000001111",
13337 => "00000010000010110000001111111111",
13338 => "00000011000001111111101000001100",
13339 => "11110101000000011111011011110101",
13340 => "00000011111110100000001011111110",
13341 => "11111010111101000000001100000100",
13342 => "00000000111110001111100011111111",
13343 => "11111110111110011111011111111001",
13344 => "11110100000000011111100000000001",
13345 => "11111001111101010000101011111101",
13346 => "11110101111111001111101100000011",
13347 => "11111100111101011111110111110110",
13348 => "11111001111111101111010111110101",
13349 => "00000100111110101111010100000000",
13350 => "00000000111111101111110111110011",
13351 => "11111000000010111111110000001010",
13352 => "11101010111111001111010111110100",
13353 => "11111001000000011110010011111100",
13354 => "11111100111111111111100111110110",
13355 => "11110011110111001111101000000000",
13356 => "11111000111100111111111000000001",
13357 => "00000010111111001110111111111110",
13358 => "11111110111110001111101111110000",
13359 => "11110100111010110000011100001001",
13360 => "11111001111110001111010011111000",
13361 => "11110011111101010000101100000001",
13362 => "00000010111111001111110111111100",
13363 => "11110110111101010000000000000010",
13364 => "11101111111010011111011100000010",
13365 => "11111011000001011110101100000011",
13366 => "11101110111100100000010111101110",
13367 => "00000101000000111110100000001011",
13368 => "11000011111111111111010011110001",
13369 => "11111100111101111111100111111100",
13370 => "00000010000001100000100111101100",
13371 => "11111011000001011111110100001100",
13372 => "11111010111110001111111011111100",
13373 => "00001000000000001111011000000110",
13374 => "11100110111111010000001111110010",
13375 => "00001000000000111101001100010011",
13376 => "11100100000000011110110111110011",
13377 => "00000010111110000000000011111010",
13378 => "11111101000001010000011011111100",
13379 => "11101101000010111110111100001101",
13380 => "11111010111011100000001111111110",
13381 => "00000100000000111111001000001000",
13382 => "11100100111111001111110111110000",
13383 => "11111110000010011101111011100110",
13384 => "11110011111111111101110111111001",
13385 => "11111101111100110000010000000100",
13386 => "00000010111110011111100011110011",
13387 => "11110011000100011111011011111101",
13388 => "11110011111111101110110011110000",
13389 => "00001100111110111110100000001110",
13390 => "11111110111101101111011000000101",
13391 => "00000011000001101110001011010101",
13392 => "00010001000001011111100011111111",
13393 => "00000100110111111101100111110011",
13394 => "11111010111111011111101111111011",
13395 => "11110000000001011111010011111010",
13396 => "11111001111111001111011111110100",
13397 => "00000011000001101111101000001010",
13398 => "00000010111110011111110100011101",
13399 => "00001000111110100000010011001110",
13400 => "00001110000000101111110000000101",
13401 => "00000110111011001111000111111110",
13402 => "11111110111101111111100000000100",
13403 => "11110111111111111111111111111101",
13404 => "11111000111111001110111011110100",
13405 => "00000100000000011111111100000000",
13406 => "11111110111111101111111100001110",
13407 => "11111101111110000000001111011000",
13408 => "00010011111111101111100100001011",
13409 => "00000000111100101110010011111011",
13410 => "11111111111101111111010000000010",
13411 => "00000000000000011111110111110111",
13412 => "11111000000001111110110011111111",
13413 => "00001001000001101111010100001000",
13414 => "11111100000001110000001000000011",
13415 => "00000100111100110000000011100101",
13416 => "00000110000001000001000100000000",
13417 => "11111010000000101111101111111111",
13418 => "11111111000001101111100111111010",
13419 => "00010000000010100000101111111011",
13420 => "11111000000001011111001000000010",
13421 => "11110111111101101111111011110111",
13422 => "11111011111110100000011100001111",
13423 => "00000000000000101111101111101101",
13424 => "00001101111111000001010000000010",
13425 => "11111001000101101111000111111101",
13426 => "00001001000001010000010000000000",
13427 => "00000011000000010000000000000011",
13428 => "00010000000100110000110100000110",
13429 => "00000011000000010001000000000011",
13430 => "00000001000001101111111000010110",
13431 => "00001111000000110001101111111001",
13432 => "00001010000001110001001100001111",
13433 => "00001111000000010001101011111111",
13434 => "11111011111111000000001100001111",
13435 => "11111101000010001111011000000010",
13436 => "00010000000010110000111111111111",
13437 => "00000111111111000000111111111101",
13438 => "11111101000011110000001011111100",
13439 => "00000000000010011111111000001101",
13440 => "00000001000001100000000100001011",
13441 => "11111100000001000000110000000001",
13442 => "11111011111111000000001100001111",
13443 => "11111000000000111111110011111110",
13444 => "11101110000000111111111100000000",
13445 => "11110101000000001110010111110100",
13446 => "11111011111110101111110011111101",
13447 => "11111100000000110000000100000100",
13448 => "00000010111100101111111111101110",
13449 => "00000001111111110000011000000000",
13450 => "11111110111111101111011011101011",
13451 => "11111101000000101111100100001111",
13452 => "00000111000010001111100000000101",
13453 => "00010001111111110000001000010000",
13454 => "11111111111111110000010000000011",
13455 => "00000001111011100000000000010110",
13456 => "11111100000011010000011100001110",
13457 => "11111110000010010001000111111111",
13458 => "11111101000010010000000100001101",
13459 => "11111110000010110000000100010101",
13460 => "11111111111110111111101000001010",
13461 => "00010010000010011111110000001110",
13462 => "11110110000011010000001111111010",
13463 => "11111011000100100001010100001010",
13464 => "00010111000001001111011111111010",
13465 => "11111101000010010010001011111101",
13466 => "00001000000010001111110111111010",
13467 => "00000010000110001111111100000101",
13468 => "00001000000001010000110100000011",
13469 => "00010001000000110000011000010010",
13470 => "00000000111111000000010011111110",
13471 => "00001010000100000001000000010010",
13472 => "00011000000011100000101000000101",
13473 => "00010110111111010001011011111010",
13474 => "00000011111110010000101100000111",
13475 => "00000100000011100000001100001101",
13476 => "00001110111110110000110100000111",
13477 => "00010001111110110000101100001011",
13478 => "00000011111111100000001100000111",
13479 => "00001000000001001110101000001010",
13480 => "00011110000010011111100000001011",
13481 => "00000101000000010000111011111001",
13482 => "00000011000000000000001000000111",
13483 => "00000011000100010000110000000001",
13484 => "00000111000010010000000011111101",
13485 => "00010011000001111111111000000001",
13486 => "11110101000001000000010011111011",
13487 => "00000011000011001111001000000110",
13488 => "00011010000010110000011000001010",
13489 => "00001101000001011111110011111010",
13490 => "00000100000000010000011100001001",
13491 => "00000010000100010000011000001010",
13492 => "00000011000001101111110000000000",
13493 => "00011001111110111111101100011010",
13494 => "00000000111101010000001100001001",
13495 => "00000010000000001110001100000100",
13496 => "00010011000011100000111000000001",
13497 => "00000000000010001111010111111101",
13498 => "00000101000010010000010100000011",
13499 => "00000100000010010000001000000011",
13500 => "00000010000100000000001100000000",
13501 => "00010100000000000000000000001101",
13502 => "11111101000000100000011111111110",
13503 => "11111110111111110000010011101110",
13504 => "00100100000001000000101111111110",
13505 => "00000111000010111111000011111110",
13506 => "00000100000010000000001111111100",
13507 => "11111010000100101111111000001100",
13508 => "00000010000010001111110100000000",
13509 => "00100001111111101111110100011100",
13510 => "11111100111111010000011100000011",
13511 => "00010010000001011111100111101010",
13512 => "00100100000100100000011100000110",
13513 => "00010101000000000000010011110111",
13514 => "00001001000001000000000100000000",
13515 => "00000011000001010000000000000101",
13516 => "00000011000010100000001000001011",
13517 => "00100110000001100000001100011100",
13518 => "11111110000000110000010000010000",
13519 => "00010110000000000000100011101000",
13520 => "00011001000111100001100000001010",
13521 => "00010010000010000000011111110110",
13522 => "00000100000011110000111100001101",
13523 => "11111101000111011111111000000010",
13524 => "00001111000001110000100000000000",
13525 => "11111011111111101111111011110101",
13526 => "00000010000100100000011111110110",
13527 => "11111011000101000000101111110101",
13528 => "00011100111111111111001000000000",
13529 => "11111111111101010000110011111011",
13530 => "00000101111111110000100000001011",
13531 => "00001111111111000001000000000010",
13532 => "00001011000011010000011011111011",
13533 => "00000011000001000000100111111001",
13534 => "11111111000000100000011000000010",
13535 => "00010010000000011111011011111111",
13536 => "11110111111111010001010100001100",
13537 => "00010101000011011111000111111110",
13538 => "00000010000001000000001000001000",
13539 => "11111101111110111111111100000100",
13540 => "11111011111111111111111100000101",
13541 => "00001100000010001111101011111110",
13542 => "00000010111111010000000111111110",
13543 => "11111101111101110000001011111100",
13544 => "11111110000001001111110000000000",
13545 => "11111011000001100001000011111111",
13546 => "00000000000000000000000111111011",
13547 => "00000000000000000000000000000000",
13548 => "00000000000000000000000000000000",
13549 => "00000000000000000000000000000000"    
);

begin

clock : process(clk)
begin
    if rising_edge(clk) then
        weights1 <= data1;
        weights2 <= data2;
        weights3 <= data3;
        weights4 <= data4;
        weights5 <= data5;
        weights6 <= data6;
        weights7 <= data7;
        weights8 <= data8;
        weights9 <= data9;
        weights10 <= data10;
    end if;
end process;

process (romAddress)
begin
    case romAddress is
        when "00000000000" => 
 data1 <= my_rom(0); 
 data2 <= my_rom(1355); 
 data3 <= my_rom(2710); 
 data4 <= my_rom(4065); 
 data5 <= my_rom(5420); 
 data6 <= my_rom(6775); 
 data7 <= my_rom(8130); 
 data8 <= my_rom(9485); 
 data9 <= my_rom(10840); 
 data10 <= my_rom(12195);
when "00000000001" => 
 data1 <= my_rom(1); 
 data2 <= my_rom(1356); 
 data3 <= my_rom(2711); 
 data4 <= my_rom(4066); 
 data5 <= my_rom(5421); 
 data6 <= my_rom(6776); 
 data7 <= my_rom(8131); 
 data8 <= my_rom(9486); 
 data9 <= my_rom(10841); 
 data10 <= my_rom(12196);
when "00000000010" => 
 data1 <= my_rom(2); 
 data2 <= my_rom(1357); 
 data3 <= my_rom(2712); 
 data4 <= my_rom(4067); 
 data5 <= my_rom(5422); 
 data6 <= my_rom(6777); 
 data7 <= my_rom(8132); 
 data8 <= my_rom(9487); 
 data9 <= my_rom(10842); 
 data10 <= my_rom(12197);
when "00000000011" => 
 data1 <= my_rom(3); 
 data2 <= my_rom(1358); 
 data3 <= my_rom(2713); 
 data4 <= my_rom(4068); 
 data5 <= my_rom(5423); 
 data6 <= my_rom(6778); 
 data7 <= my_rom(8133); 
 data8 <= my_rom(9488); 
 data9 <= my_rom(10843); 
 data10 <= my_rom(12198);
when "00000000100" => 
 data1 <= my_rom(4); 
 data2 <= my_rom(1359); 
 data3 <= my_rom(2714); 
 data4 <= my_rom(4069); 
 data5 <= my_rom(5424); 
 data6 <= my_rom(6779); 
 data7 <= my_rom(8134); 
 data8 <= my_rom(9489); 
 data9 <= my_rom(10844); 
 data10 <= my_rom(12199);
when "00000000101" => 
 data1 <= my_rom(5); 
 data2 <= my_rom(1360); 
 data3 <= my_rom(2715); 
 data4 <= my_rom(4070); 
 data5 <= my_rom(5425); 
 data6 <= my_rom(6780); 
 data7 <= my_rom(8135); 
 data8 <= my_rom(9490); 
 data9 <= my_rom(10845); 
 data10 <= my_rom(12200);
when "00000000110" => 
 data1 <= my_rom(6); 
 data2 <= my_rom(1361); 
 data3 <= my_rom(2716); 
 data4 <= my_rom(4071); 
 data5 <= my_rom(5426); 
 data6 <= my_rom(6781); 
 data7 <= my_rom(8136); 
 data8 <= my_rom(9491); 
 data9 <= my_rom(10846); 
 data10 <= my_rom(12201);
when "00000000111" => 
 data1 <= my_rom(7); 
 data2 <= my_rom(1362); 
 data3 <= my_rom(2717); 
 data4 <= my_rom(4072); 
 data5 <= my_rom(5427); 
 data6 <= my_rom(6782); 
 data7 <= my_rom(8137); 
 data8 <= my_rom(9492); 
 data9 <= my_rom(10847); 
 data10 <= my_rom(12202);
when "00000001000" => 
 data1 <= my_rom(8); 
 data2 <= my_rom(1363); 
 data3 <= my_rom(2718); 
 data4 <= my_rom(4073); 
 data5 <= my_rom(5428); 
 data6 <= my_rom(6783); 
 data7 <= my_rom(8138); 
 data8 <= my_rom(9493); 
 data9 <= my_rom(10848); 
 data10 <= my_rom(12203);
when "00000001001" => 
 data1 <= my_rom(9); 
 data2 <= my_rom(1364); 
 data3 <= my_rom(2719); 
 data4 <= my_rom(4074); 
 data5 <= my_rom(5429); 
 data6 <= my_rom(6784); 
 data7 <= my_rom(8139); 
 data8 <= my_rom(9494); 
 data9 <= my_rom(10849); 
 data10 <= my_rom(12204);
when "00000001010" => 
 data1 <= my_rom(10); 
 data2 <= my_rom(1365); 
 data3 <= my_rom(2720); 
 data4 <= my_rom(4075); 
 data5 <= my_rom(5430); 
 data6 <= my_rom(6785); 
 data7 <= my_rom(8140); 
 data8 <= my_rom(9495); 
 data9 <= my_rom(10850); 
 data10 <= my_rom(12205);
when "00000001011" => 
 data1 <= my_rom(11); 
 data2 <= my_rom(1366); 
 data3 <= my_rom(2721); 
 data4 <= my_rom(4076); 
 data5 <= my_rom(5431); 
 data6 <= my_rom(6786); 
 data7 <= my_rom(8141); 
 data8 <= my_rom(9496); 
 data9 <= my_rom(10851); 
 data10 <= my_rom(12206);
when "00000001100" => 
 data1 <= my_rom(12); 
 data2 <= my_rom(1367); 
 data3 <= my_rom(2722); 
 data4 <= my_rom(4077); 
 data5 <= my_rom(5432); 
 data6 <= my_rom(6787); 
 data7 <= my_rom(8142); 
 data8 <= my_rom(9497); 
 data9 <= my_rom(10852); 
 data10 <= my_rom(12207);
when "00000001101" => 
 data1 <= my_rom(13); 
 data2 <= my_rom(1368); 
 data3 <= my_rom(2723); 
 data4 <= my_rom(4078); 
 data5 <= my_rom(5433); 
 data6 <= my_rom(6788); 
 data7 <= my_rom(8143); 
 data8 <= my_rom(9498); 
 data9 <= my_rom(10853); 
 data10 <= my_rom(12208);
when "00000001110" => 
 data1 <= my_rom(14); 
 data2 <= my_rom(1369); 
 data3 <= my_rom(2724); 
 data4 <= my_rom(4079); 
 data5 <= my_rom(5434); 
 data6 <= my_rom(6789); 
 data7 <= my_rom(8144); 
 data8 <= my_rom(9499); 
 data9 <= my_rom(10854); 
 data10 <= my_rom(12209);
when "00000001111" => 
 data1 <= my_rom(15); 
 data2 <= my_rom(1370); 
 data3 <= my_rom(2725); 
 data4 <= my_rom(4080); 
 data5 <= my_rom(5435); 
 data6 <= my_rom(6790); 
 data7 <= my_rom(8145); 
 data8 <= my_rom(9500); 
 data9 <= my_rom(10855); 
 data10 <= my_rom(12210);
when "00000010000" => 
 data1 <= my_rom(16); 
 data2 <= my_rom(1371); 
 data3 <= my_rom(2726); 
 data4 <= my_rom(4081); 
 data5 <= my_rom(5436); 
 data6 <= my_rom(6791); 
 data7 <= my_rom(8146); 
 data8 <= my_rom(9501); 
 data9 <= my_rom(10856); 
 data10 <= my_rom(12211);
when "00000010001" => 
 data1 <= my_rom(17); 
 data2 <= my_rom(1372); 
 data3 <= my_rom(2727); 
 data4 <= my_rom(4082); 
 data5 <= my_rom(5437); 
 data6 <= my_rom(6792); 
 data7 <= my_rom(8147); 
 data8 <= my_rom(9502); 
 data9 <= my_rom(10857); 
 data10 <= my_rom(12212);
when "00000010010" => 
 data1 <= my_rom(18); 
 data2 <= my_rom(1373); 
 data3 <= my_rom(2728); 
 data4 <= my_rom(4083); 
 data5 <= my_rom(5438); 
 data6 <= my_rom(6793); 
 data7 <= my_rom(8148); 
 data8 <= my_rom(9503); 
 data9 <= my_rom(10858); 
 data10 <= my_rom(12213);
when "00000010011" => 
 data1 <= my_rom(19); 
 data2 <= my_rom(1374); 
 data3 <= my_rom(2729); 
 data4 <= my_rom(4084); 
 data5 <= my_rom(5439); 
 data6 <= my_rom(6794); 
 data7 <= my_rom(8149); 
 data8 <= my_rom(9504); 
 data9 <= my_rom(10859); 
 data10 <= my_rom(12214);
when "00000010100" => 
 data1 <= my_rom(20); 
 data2 <= my_rom(1375); 
 data3 <= my_rom(2730); 
 data4 <= my_rom(4085); 
 data5 <= my_rom(5440); 
 data6 <= my_rom(6795); 
 data7 <= my_rom(8150); 
 data8 <= my_rom(9505); 
 data9 <= my_rom(10860); 
 data10 <= my_rom(12215);
when "00000010101" => 
 data1 <= my_rom(21); 
 data2 <= my_rom(1376); 
 data3 <= my_rom(2731); 
 data4 <= my_rom(4086); 
 data5 <= my_rom(5441); 
 data6 <= my_rom(6796); 
 data7 <= my_rom(8151); 
 data8 <= my_rom(9506); 
 data9 <= my_rom(10861); 
 data10 <= my_rom(12216);
when "00000010110" => 
 data1 <= my_rom(22); 
 data2 <= my_rom(1377); 
 data3 <= my_rom(2732); 
 data4 <= my_rom(4087); 
 data5 <= my_rom(5442); 
 data6 <= my_rom(6797); 
 data7 <= my_rom(8152); 
 data8 <= my_rom(9507); 
 data9 <= my_rom(10862); 
 data10 <= my_rom(12217);
when "00000010111" => 
 data1 <= my_rom(23); 
 data2 <= my_rom(1378); 
 data3 <= my_rom(2733); 
 data4 <= my_rom(4088); 
 data5 <= my_rom(5443); 
 data6 <= my_rom(6798); 
 data7 <= my_rom(8153); 
 data8 <= my_rom(9508); 
 data9 <= my_rom(10863); 
 data10 <= my_rom(12218);
when "00000011000" => 
 data1 <= my_rom(24); 
 data2 <= my_rom(1379); 
 data3 <= my_rom(2734); 
 data4 <= my_rom(4089); 
 data5 <= my_rom(5444); 
 data6 <= my_rom(6799); 
 data7 <= my_rom(8154); 
 data8 <= my_rom(9509); 
 data9 <= my_rom(10864); 
 data10 <= my_rom(12219);
when "00000011001" => 
 data1 <= my_rom(25); 
 data2 <= my_rom(1380); 
 data3 <= my_rom(2735); 
 data4 <= my_rom(4090); 
 data5 <= my_rom(5445); 
 data6 <= my_rom(6800); 
 data7 <= my_rom(8155); 
 data8 <= my_rom(9510); 
 data9 <= my_rom(10865); 
 data10 <= my_rom(12220);
when "00000011010" => 
 data1 <= my_rom(26); 
 data2 <= my_rom(1381); 
 data3 <= my_rom(2736); 
 data4 <= my_rom(4091); 
 data5 <= my_rom(5446); 
 data6 <= my_rom(6801); 
 data7 <= my_rom(8156); 
 data8 <= my_rom(9511); 
 data9 <= my_rom(10866); 
 data10 <= my_rom(12221);
when "00000011011" => 
 data1 <= my_rom(27); 
 data2 <= my_rom(1382); 
 data3 <= my_rom(2737); 
 data4 <= my_rom(4092); 
 data5 <= my_rom(5447); 
 data6 <= my_rom(6802); 
 data7 <= my_rom(8157); 
 data8 <= my_rom(9512); 
 data9 <= my_rom(10867); 
 data10 <= my_rom(12222);
when "00000011100" => 
 data1 <= my_rom(28); 
 data2 <= my_rom(1383); 
 data3 <= my_rom(2738); 
 data4 <= my_rom(4093); 
 data5 <= my_rom(5448); 
 data6 <= my_rom(6803); 
 data7 <= my_rom(8158); 
 data8 <= my_rom(9513); 
 data9 <= my_rom(10868); 
 data10 <= my_rom(12223);
when "00000011101" => 
 data1 <= my_rom(29); 
 data2 <= my_rom(1384); 
 data3 <= my_rom(2739); 
 data4 <= my_rom(4094); 
 data5 <= my_rom(5449); 
 data6 <= my_rom(6804); 
 data7 <= my_rom(8159); 
 data8 <= my_rom(9514); 
 data9 <= my_rom(10869); 
 data10 <= my_rom(12224);
when "00000011110" => 
 data1 <= my_rom(30); 
 data2 <= my_rom(1385); 
 data3 <= my_rom(2740); 
 data4 <= my_rom(4095); 
 data5 <= my_rom(5450); 
 data6 <= my_rom(6805); 
 data7 <= my_rom(8160); 
 data8 <= my_rom(9515); 
 data9 <= my_rom(10870); 
 data10 <= my_rom(12225);
when "00000011111" => 
 data1 <= my_rom(31); 
 data2 <= my_rom(1386); 
 data3 <= my_rom(2741); 
 data4 <= my_rom(4096); 
 data5 <= my_rom(5451); 
 data6 <= my_rom(6806); 
 data7 <= my_rom(8161); 
 data8 <= my_rom(9516); 
 data9 <= my_rom(10871); 
 data10 <= my_rom(12226);
when "00000100000" => 
 data1 <= my_rom(32); 
 data2 <= my_rom(1387); 
 data3 <= my_rom(2742); 
 data4 <= my_rom(4097); 
 data5 <= my_rom(5452); 
 data6 <= my_rom(6807); 
 data7 <= my_rom(8162); 
 data8 <= my_rom(9517); 
 data9 <= my_rom(10872); 
 data10 <= my_rom(12227);
when "00000100001" => 
 data1 <= my_rom(33); 
 data2 <= my_rom(1388); 
 data3 <= my_rom(2743); 
 data4 <= my_rom(4098); 
 data5 <= my_rom(5453); 
 data6 <= my_rom(6808); 
 data7 <= my_rom(8163); 
 data8 <= my_rom(9518); 
 data9 <= my_rom(10873); 
 data10 <= my_rom(12228);
when "00000100010" => 
 data1 <= my_rom(34); 
 data2 <= my_rom(1389); 
 data3 <= my_rom(2744); 
 data4 <= my_rom(4099); 
 data5 <= my_rom(5454); 
 data6 <= my_rom(6809); 
 data7 <= my_rom(8164); 
 data8 <= my_rom(9519); 
 data9 <= my_rom(10874); 
 data10 <= my_rom(12229);
when "00000100011" => 
 data1 <= my_rom(35); 
 data2 <= my_rom(1390); 
 data3 <= my_rom(2745); 
 data4 <= my_rom(4100); 
 data5 <= my_rom(5455); 
 data6 <= my_rom(6810); 
 data7 <= my_rom(8165); 
 data8 <= my_rom(9520); 
 data9 <= my_rom(10875); 
 data10 <= my_rom(12230);
when "00000100100" => 
 data1 <= my_rom(36); 
 data2 <= my_rom(1391); 
 data3 <= my_rom(2746); 
 data4 <= my_rom(4101); 
 data5 <= my_rom(5456); 
 data6 <= my_rom(6811); 
 data7 <= my_rom(8166); 
 data8 <= my_rom(9521); 
 data9 <= my_rom(10876); 
 data10 <= my_rom(12231);
when "00000100101" => 
 data1 <= my_rom(37); 
 data2 <= my_rom(1392); 
 data3 <= my_rom(2747); 
 data4 <= my_rom(4102); 
 data5 <= my_rom(5457); 
 data6 <= my_rom(6812); 
 data7 <= my_rom(8167); 
 data8 <= my_rom(9522); 
 data9 <= my_rom(10877); 
 data10 <= my_rom(12232);
when "00000100110" => 
 data1 <= my_rom(38); 
 data2 <= my_rom(1393); 
 data3 <= my_rom(2748); 
 data4 <= my_rom(4103); 
 data5 <= my_rom(5458); 
 data6 <= my_rom(6813); 
 data7 <= my_rom(8168); 
 data8 <= my_rom(9523); 
 data9 <= my_rom(10878); 
 data10 <= my_rom(12233);
when "00000100111" => 
 data1 <= my_rom(39); 
 data2 <= my_rom(1394); 
 data3 <= my_rom(2749); 
 data4 <= my_rom(4104); 
 data5 <= my_rom(5459); 
 data6 <= my_rom(6814); 
 data7 <= my_rom(8169); 
 data8 <= my_rom(9524); 
 data9 <= my_rom(10879); 
 data10 <= my_rom(12234);
when "00000101000" => 
 data1 <= my_rom(40); 
 data2 <= my_rom(1395); 
 data3 <= my_rom(2750); 
 data4 <= my_rom(4105); 
 data5 <= my_rom(5460); 
 data6 <= my_rom(6815); 
 data7 <= my_rom(8170); 
 data8 <= my_rom(9525); 
 data9 <= my_rom(10880); 
 data10 <= my_rom(12235);
when "00000101001" => 
 data1 <= my_rom(41); 
 data2 <= my_rom(1396); 
 data3 <= my_rom(2751); 
 data4 <= my_rom(4106); 
 data5 <= my_rom(5461); 
 data6 <= my_rom(6816); 
 data7 <= my_rom(8171); 
 data8 <= my_rom(9526); 
 data9 <= my_rom(10881); 
 data10 <= my_rom(12236);
when "00000101010" => 
 data1 <= my_rom(42); 
 data2 <= my_rom(1397); 
 data3 <= my_rom(2752); 
 data4 <= my_rom(4107); 
 data5 <= my_rom(5462); 
 data6 <= my_rom(6817); 
 data7 <= my_rom(8172); 
 data8 <= my_rom(9527); 
 data9 <= my_rom(10882); 
 data10 <= my_rom(12237);
when "00000101011" => 
 data1 <= my_rom(43); 
 data2 <= my_rom(1398); 
 data3 <= my_rom(2753); 
 data4 <= my_rom(4108); 
 data5 <= my_rom(5463); 
 data6 <= my_rom(6818); 
 data7 <= my_rom(8173); 
 data8 <= my_rom(9528); 
 data9 <= my_rom(10883); 
 data10 <= my_rom(12238);
when "00000101100" => 
 data1 <= my_rom(44); 
 data2 <= my_rom(1399); 
 data3 <= my_rom(2754); 
 data4 <= my_rom(4109); 
 data5 <= my_rom(5464); 
 data6 <= my_rom(6819); 
 data7 <= my_rom(8174); 
 data8 <= my_rom(9529); 
 data9 <= my_rom(10884); 
 data10 <= my_rom(12239);
when "00000101101" => 
 data1 <= my_rom(45); 
 data2 <= my_rom(1400); 
 data3 <= my_rom(2755); 
 data4 <= my_rom(4110); 
 data5 <= my_rom(5465); 
 data6 <= my_rom(6820); 
 data7 <= my_rom(8175); 
 data8 <= my_rom(9530); 
 data9 <= my_rom(10885); 
 data10 <= my_rom(12240);
when "00000101110" => 
 data1 <= my_rom(46); 
 data2 <= my_rom(1401); 
 data3 <= my_rom(2756); 
 data4 <= my_rom(4111); 
 data5 <= my_rom(5466); 
 data6 <= my_rom(6821); 
 data7 <= my_rom(8176); 
 data8 <= my_rom(9531); 
 data9 <= my_rom(10886); 
 data10 <= my_rom(12241);
when "00000101111" => 
 data1 <= my_rom(47); 
 data2 <= my_rom(1402); 
 data3 <= my_rom(2757); 
 data4 <= my_rom(4112); 
 data5 <= my_rom(5467); 
 data6 <= my_rom(6822); 
 data7 <= my_rom(8177); 
 data8 <= my_rom(9532); 
 data9 <= my_rom(10887); 
 data10 <= my_rom(12242);
when "00000110000" => 
 data1 <= my_rom(48); 
 data2 <= my_rom(1403); 
 data3 <= my_rom(2758); 
 data4 <= my_rom(4113); 
 data5 <= my_rom(5468); 
 data6 <= my_rom(6823); 
 data7 <= my_rom(8178); 
 data8 <= my_rom(9533); 
 data9 <= my_rom(10888); 
 data10 <= my_rom(12243);
when "00000110001" => 
 data1 <= my_rom(49); 
 data2 <= my_rom(1404); 
 data3 <= my_rom(2759); 
 data4 <= my_rom(4114); 
 data5 <= my_rom(5469); 
 data6 <= my_rom(6824); 
 data7 <= my_rom(8179); 
 data8 <= my_rom(9534); 
 data9 <= my_rom(10889); 
 data10 <= my_rom(12244);
when "00000110010" => 
 data1 <= my_rom(50); 
 data2 <= my_rom(1405); 
 data3 <= my_rom(2760); 
 data4 <= my_rom(4115); 
 data5 <= my_rom(5470); 
 data6 <= my_rom(6825); 
 data7 <= my_rom(8180); 
 data8 <= my_rom(9535); 
 data9 <= my_rom(10890); 
 data10 <= my_rom(12245);
when "00000110011" => 
 data1 <= my_rom(51); 
 data2 <= my_rom(1406); 
 data3 <= my_rom(2761); 
 data4 <= my_rom(4116); 
 data5 <= my_rom(5471); 
 data6 <= my_rom(6826); 
 data7 <= my_rom(8181); 
 data8 <= my_rom(9536); 
 data9 <= my_rom(10891); 
 data10 <= my_rom(12246);
when "00000110100" => 
 data1 <= my_rom(52); 
 data2 <= my_rom(1407); 
 data3 <= my_rom(2762); 
 data4 <= my_rom(4117); 
 data5 <= my_rom(5472); 
 data6 <= my_rom(6827); 
 data7 <= my_rom(8182); 
 data8 <= my_rom(9537); 
 data9 <= my_rom(10892); 
 data10 <= my_rom(12247);
when "00000110101" => 
 data1 <= my_rom(53); 
 data2 <= my_rom(1408); 
 data3 <= my_rom(2763); 
 data4 <= my_rom(4118); 
 data5 <= my_rom(5473); 
 data6 <= my_rom(6828); 
 data7 <= my_rom(8183); 
 data8 <= my_rom(9538); 
 data9 <= my_rom(10893); 
 data10 <= my_rom(12248);
when "00000110110" => 
 data1 <= my_rom(54); 
 data2 <= my_rom(1409); 
 data3 <= my_rom(2764); 
 data4 <= my_rom(4119); 
 data5 <= my_rom(5474); 
 data6 <= my_rom(6829); 
 data7 <= my_rom(8184); 
 data8 <= my_rom(9539); 
 data9 <= my_rom(10894); 
 data10 <= my_rom(12249);
when "00000110111" => 
 data1 <= my_rom(55); 
 data2 <= my_rom(1410); 
 data3 <= my_rom(2765); 
 data4 <= my_rom(4120); 
 data5 <= my_rom(5475); 
 data6 <= my_rom(6830); 
 data7 <= my_rom(8185); 
 data8 <= my_rom(9540); 
 data9 <= my_rom(10895); 
 data10 <= my_rom(12250);
when "00000111000" => 
 data1 <= my_rom(56); 
 data2 <= my_rom(1411); 
 data3 <= my_rom(2766); 
 data4 <= my_rom(4121); 
 data5 <= my_rom(5476); 
 data6 <= my_rom(6831); 
 data7 <= my_rom(8186); 
 data8 <= my_rom(9541); 
 data9 <= my_rom(10896); 
 data10 <= my_rom(12251);
when "00000111001" => 
 data1 <= my_rom(57); 
 data2 <= my_rom(1412); 
 data3 <= my_rom(2767); 
 data4 <= my_rom(4122); 
 data5 <= my_rom(5477); 
 data6 <= my_rom(6832); 
 data7 <= my_rom(8187); 
 data8 <= my_rom(9542); 
 data9 <= my_rom(10897); 
 data10 <= my_rom(12252);
when "00000111010" => 
 data1 <= my_rom(58); 
 data2 <= my_rom(1413); 
 data3 <= my_rom(2768); 
 data4 <= my_rom(4123); 
 data5 <= my_rom(5478); 
 data6 <= my_rom(6833); 
 data7 <= my_rom(8188); 
 data8 <= my_rom(9543); 
 data9 <= my_rom(10898); 
 data10 <= my_rom(12253);
when "00000111011" => 
 data1 <= my_rom(59); 
 data2 <= my_rom(1414); 
 data3 <= my_rom(2769); 
 data4 <= my_rom(4124); 
 data5 <= my_rom(5479); 
 data6 <= my_rom(6834); 
 data7 <= my_rom(8189); 
 data8 <= my_rom(9544); 
 data9 <= my_rom(10899); 
 data10 <= my_rom(12254);
when "00000111100" => 
 data1 <= my_rom(60); 
 data2 <= my_rom(1415); 
 data3 <= my_rom(2770); 
 data4 <= my_rom(4125); 
 data5 <= my_rom(5480); 
 data6 <= my_rom(6835); 
 data7 <= my_rom(8190); 
 data8 <= my_rom(9545); 
 data9 <= my_rom(10900); 
 data10 <= my_rom(12255);
when "00000111101" => 
 data1 <= my_rom(61); 
 data2 <= my_rom(1416); 
 data3 <= my_rom(2771); 
 data4 <= my_rom(4126); 
 data5 <= my_rom(5481); 
 data6 <= my_rom(6836); 
 data7 <= my_rom(8191); 
 data8 <= my_rom(9546); 
 data9 <= my_rom(10901); 
 data10 <= my_rom(12256);
when "00000111110" => 
 data1 <= my_rom(62); 
 data2 <= my_rom(1417); 
 data3 <= my_rom(2772); 
 data4 <= my_rom(4127); 
 data5 <= my_rom(5482); 
 data6 <= my_rom(6837); 
 data7 <= my_rom(8192); 
 data8 <= my_rom(9547); 
 data9 <= my_rom(10902); 
 data10 <= my_rom(12257);
when "00000111111" => 
 data1 <= my_rom(63); 
 data2 <= my_rom(1418); 
 data3 <= my_rom(2773); 
 data4 <= my_rom(4128); 
 data5 <= my_rom(5483); 
 data6 <= my_rom(6838); 
 data7 <= my_rom(8193); 
 data8 <= my_rom(9548); 
 data9 <= my_rom(10903); 
 data10 <= my_rom(12258);
when "00001000000" => 
 data1 <= my_rom(64); 
 data2 <= my_rom(1419); 
 data3 <= my_rom(2774); 
 data4 <= my_rom(4129); 
 data5 <= my_rom(5484); 
 data6 <= my_rom(6839); 
 data7 <= my_rom(8194); 
 data8 <= my_rom(9549); 
 data9 <= my_rom(10904); 
 data10 <= my_rom(12259);
when "00001000001" => 
 data1 <= my_rom(65); 
 data2 <= my_rom(1420); 
 data3 <= my_rom(2775); 
 data4 <= my_rom(4130); 
 data5 <= my_rom(5485); 
 data6 <= my_rom(6840); 
 data7 <= my_rom(8195); 
 data8 <= my_rom(9550); 
 data9 <= my_rom(10905); 
 data10 <= my_rom(12260);
when "00001000010" => 
 data1 <= my_rom(66); 
 data2 <= my_rom(1421); 
 data3 <= my_rom(2776); 
 data4 <= my_rom(4131); 
 data5 <= my_rom(5486); 
 data6 <= my_rom(6841); 
 data7 <= my_rom(8196); 
 data8 <= my_rom(9551); 
 data9 <= my_rom(10906); 
 data10 <= my_rom(12261);
when "00001000011" => 
 data1 <= my_rom(67); 
 data2 <= my_rom(1422); 
 data3 <= my_rom(2777); 
 data4 <= my_rom(4132); 
 data5 <= my_rom(5487); 
 data6 <= my_rom(6842); 
 data7 <= my_rom(8197); 
 data8 <= my_rom(9552); 
 data9 <= my_rom(10907); 
 data10 <= my_rom(12262);
when "00001000100" => 
 data1 <= my_rom(68); 
 data2 <= my_rom(1423); 
 data3 <= my_rom(2778); 
 data4 <= my_rom(4133); 
 data5 <= my_rom(5488); 
 data6 <= my_rom(6843); 
 data7 <= my_rom(8198); 
 data8 <= my_rom(9553); 
 data9 <= my_rom(10908); 
 data10 <= my_rom(12263);
when "00001000101" => 
 data1 <= my_rom(69); 
 data2 <= my_rom(1424); 
 data3 <= my_rom(2779); 
 data4 <= my_rom(4134); 
 data5 <= my_rom(5489); 
 data6 <= my_rom(6844); 
 data7 <= my_rom(8199); 
 data8 <= my_rom(9554); 
 data9 <= my_rom(10909); 
 data10 <= my_rom(12264);
when "00001000110" => 
 data1 <= my_rom(70); 
 data2 <= my_rom(1425); 
 data3 <= my_rom(2780); 
 data4 <= my_rom(4135); 
 data5 <= my_rom(5490); 
 data6 <= my_rom(6845); 
 data7 <= my_rom(8200); 
 data8 <= my_rom(9555); 
 data9 <= my_rom(10910); 
 data10 <= my_rom(12265);
when "00001000111" => 
 data1 <= my_rom(71); 
 data2 <= my_rom(1426); 
 data3 <= my_rom(2781); 
 data4 <= my_rom(4136); 
 data5 <= my_rom(5491); 
 data6 <= my_rom(6846); 
 data7 <= my_rom(8201); 
 data8 <= my_rom(9556); 
 data9 <= my_rom(10911); 
 data10 <= my_rom(12266);
when "00001001000" => 
 data1 <= my_rom(72); 
 data2 <= my_rom(1427); 
 data3 <= my_rom(2782); 
 data4 <= my_rom(4137); 
 data5 <= my_rom(5492); 
 data6 <= my_rom(6847); 
 data7 <= my_rom(8202); 
 data8 <= my_rom(9557); 
 data9 <= my_rom(10912); 
 data10 <= my_rom(12267);
when "00001001001" => 
 data1 <= my_rom(73); 
 data2 <= my_rom(1428); 
 data3 <= my_rom(2783); 
 data4 <= my_rom(4138); 
 data5 <= my_rom(5493); 
 data6 <= my_rom(6848); 
 data7 <= my_rom(8203); 
 data8 <= my_rom(9558); 
 data9 <= my_rom(10913); 
 data10 <= my_rom(12268);
when "00001001010" => 
 data1 <= my_rom(74); 
 data2 <= my_rom(1429); 
 data3 <= my_rom(2784); 
 data4 <= my_rom(4139); 
 data5 <= my_rom(5494); 
 data6 <= my_rom(6849); 
 data7 <= my_rom(8204); 
 data8 <= my_rom(9559); 
 data9 <= my_rom(10914); 
 data10 <= my_rom(12269);
when "00001001011" => 
 data1 <= my_rom(75); 
 data2 <= my_rom(1430); 
 data3 <= my_rom(2785); 
 data4 <= my_rom(4140); 
 data5 <= my_rom(5495); 
 data6 <= my_rom(6850); 
 data7 <= my_rom(8205); 
 data8 <= my_rom(9560); 
 data9 <= my_rom(10915); 
 data10 <= my_rom(12270);
when "00001001100" => 
 data1 <= my_rom(76); 
 data2 <= my_rom(1431); 
 data3 <= my_rom(2786); 
 data4 <= my_rom(4141); 
 data5 <= my_rom(5496); 
 data6 <= my_rom(6851); 
 data7 <= my_rom(8206); 
 data8 <= my_rom(9561); 
 data9 <= my_rom(10916); 
 data10 <= my_rom(12271);
when "00001001101" => 
 data1 <= my_rom(77); 
 data2 <= my_rom(1432); 
 data3 <= my_rom(2787); 
 data4 <= my_rom(4142); 
 data5 <= my_rom(5497); 
 data6 <= my_rom(6852); 
 data7 <= my_rom(8207); 
 data8 <= my_rom(9562); 
 data9 <= my_rom(10917); 
 data10 <= my_rom(12272);
when "00001001110" => 
 data1 <= my_rom(78); 
 data2 <= my_rom(1433); 
 data3 <= my_rom(2788); 
 data4 <= my_rom(4143); 
 data5 <= my_rom(5498); 
 data6 <= my_rom(6853); 
 data7 <= my_rom(8208); 
 data8 <= my_rom(9563); 
 data9 <= my_rom(10918); 
 data10 <= my_rom(12273);
when "00001001111" => 
 data1 <= my_rom(79); 
 data2 <= my_rom(1434); 
 data3 <= my_rom(2789); 
 data4 <= my_rom(4144); 
 data5 <= my_rom(5499); 
 data6 <= my_rom(6854); 
 data7 <= my_rom(8209); 
 data8 <= my_rom(9564); 
 data9 <= my_rom(10919); 
 data10 <= my_rom(12274);
when "00001010000" => 
 data1 <= my_rom(80); 
 data2 <= my_rom(1435); 
 data3 <= my_rom(2790); 
 data4 <= my_rom(4145); 
 data5 <= my_rom(5500); 
 data6 <= my_rom(6855); 
 data7 <= my_rom(8210); 
 data8 <= my_rom(9565); 
 data9 <= my_rom(10920); 
 data10 <= my_rom(12275);
when "00001010001" => 
 data1 <= my_rom(81); 
 data2 <= my_rom(1436); 
 data3 <= my_rom(2791); 
 data4 <= my_rom(4146); 
 data5 <= my_rom(5501); 
 data6 <= my_rom(6856); 
 data7 <= my_rom(8211); 
 data8 <= my_rom(9566); 
 data9 <= my_rom(10921); 
 data10 <= my_rom(12276);
when "00001010010" => 
 data1 <= my_rom(82); 
 data2 <= my_rom(1437); 
 data3 <= my_rom(2792); 
 data4 <= my_rom(4147); 
 data5 <= my_rom(5502); 
 data6 <= my_rom(6857); 
 data7 <= my_rom(8212); 
 data8 <= my_rom(9567); 
 data9 <= my_rom(10922); 
 data10 <= my_rom(12277);
when "00001010011" => 
 data1 <= my_rom(83); 
 data2 <= my_rom(1438); 
 data3 <= my_rom(2793); 
 data4 <= my_rom(4148); 
 data5 <= my_rom(5503); 
 data6 <= my_rom(6858); 
 data7 <= my_rom(8213); 
 data8 <= my_rom(9568); 
 data9 <= my_rom(10923); 
 data10 <= my_rom(12278);
when "00001010100" => 
 data1 <= my_rom(84); 
 data2 <= my_rom(1439); 
 data3 <= my_rom(2794); 
 data4 <= my_rom(4149); 
 data5 <= my_rom(5504); 
 data6 <= my_rom(6859); 
 data7 <= my_rom(8214); 
 data8 <= my_rom(9569); 
 data9 <= my_rom(10924); 
 data10 <= my_rom(12279);
when "00001010101" => 
 data1 <= my_rom(85); 
 data2 <= my_rom(1440); 
 data3 <= my_rom(2795); 
 data4 <= my_rom(4150); 
 data5 <= my_rom(5505); 
 data6 <= my_rom(6860); 
 data7 <= my_rom(8215); 
 data8 <= my_rom(9570); 
 data9 <= my_rom(10925); 
 data10 <= my_rom(12280);
when "00001010110" => 
 data1 <= my_rom(86); 
 data2 <= my_rom(1441); 
 data3 <= my_rom(2796); 
 data4 <= my_rom(4151); 
 data5 <= my_rom(5506); 
 data6 <= my_rom(6861); 
 data7 <= my_rom(8216); 
 data8 <= my_rom(9571); 
 data9 <= my_rom(10926); 
 data10 <= my_rom(12281);
when "00001010111" => 
 data1 <= my_rom(87); 
 data2 <= my_rom(1442); 
 data3 <= my_rom(2797); 
 data4 <= my_rom(4152); 
 data5 <= my_rom(5507); 
 data6 <= my_rom(6862); 
 data7 <= my_rom(8217); 
 data8 <= my_rom(9572); 
 data9 <= my_rom(10927); 
 data10 <= my_rom(12282);
when "00001011000" => 
 data1 <= my_rom(88); 
 data2 <= my_rom(1443); 
 data3 <= my_rom(2798); 
 data4 <= my_rom(4153); 
 data5 <= my_rom(5508); 
 data6 <= my_rom(6863); 
 data7 <= my_rom(8218); 
 data8 <= my_rom(9573); 
 data9 <= my_rom(10928); 
 data10 <= my_rom(12283);
when "00001011001" => 
 data1 <= my_rom(89); 
 data2 <= my_rom(1444); 
 data3 <= my_rom(2799); 
 data4 <= my_rom(4154); 
 data5 <= my_rom(5509); 
 data6 <= my_rom(6864); 
 data7 <= my_rom(8219); 
 data8 <= my_rom(9574); 
 data9 <= my_rom(10929); 
 data10 <= my_rom(12284);
when "00001011010" => 
 data1 <= my_rom(90); 
 data2 <= my_rom(1445); 
 data3 <= my_rom(2800); 
 data4 <= my_rom(4155); 
 data5 <= my_rom(5510); 
 data6 <= my_rom(6865); 
 data7 <= my_rom(8220); 
 data8 <= my_rom(9575); 
 data9 <= my_rom(10930); 
 data10 <= my_rom(12285);
when "00001011011" => 
 data1 <= my_rom(91); 
 data2 <= my_rom(1446); 
 data3 <= my_rom(2801); 
 data4 <= my_rom(4156); 
 data5 <= my_rom(5511); 
 data6 <= my_rom(6866); 
 data7 <= my_rom(8221); 
 data8 <= my_rom(9576); 
 data9 <= my_rom(10931); 
 data10 <= my_rom(12286);
when "00001011100" => 
 data1 <= my_rom(92); 
 data2 <= my_rom(1447); 
 data3 <= my_rom(2802); 
 data4 <= my_rom(4157); 
 data5 <= my_rom(5512); 
 data6 <= my_rom(6867); 
 data7 <= my_rom(8222); 
 data8 <= my_rom(9577); 
 data9 <= my_rom(10932); 
 data10 <= my_rom(12287);
when "00001011101" => 
 data1 <= my_rom(93); 
 data2 <= my_rom(1448); 
 data3 <= my_rom(2803); 
 data4 <= my_rom(4158); 
 data5 <= my_rom(5513); 
 data6 <= my_rom(6868); 
 data7 <= my_rom(8223); 
 data8 <= my_rom(9578); 
 data9 <= my_rom(10933); 
 data10 <= my_rom(12288);
when "00001011110" => 
 data1 <= my_rom(94); 
 data2 <= my_rom(1449); 
 data3 <= my_rom(2804); 
 data4 <= my_rom(4159); 
 data5 <= my_rom(5514); 
 data6 <= my_rom(6869); 
 data7 <= my_rom(8224); 
 data8 <= my_rom(9579); 
 data9 <= my_rom(10934); 
 data10 <= my_rom(12289);
when "00001011111" => 
 data1 <= my_rom(95); 
 data2 <= my_rom(1450); 
 data3 <= my_rom(2805); 
 data4 <= my_rom(4160); 
 data5 <= my_rom(5515); 
 data6 <= my_rom(6870); 
 data7 <= my_rom(8225); 
 data8 <= my_rom(9580); 
 data9 <= my_rom(10935); 
 data10 <= my_rom(12290);
when "00001100000" => 
 data1 <= my_rom(96); 
 data2 <= my_rom(1451); 
 data3 <= my_rom(2806); 
 data4 <= my_rom(4161); 
 data5 <= my_rom(5516); 
 data6 <= my_rom(6871); 
 data7 <= my_rom(8226); 
 data8 <= my_rom(9581); 
 data9 <= my_rom(10936); 
 data10 <= my_rom(12291);
when "00001100001" => 
 data1 <= my_rom(97); 
 data2 <= my_rom(1452); 
 data3 <= my_rom(2807); 
 data4 <= my_rom(4162); 
 data5 <= my_rom(5517); 
 data6 <= my_rom(6872); 
 data7 <= my_rom(8227); 
 data8 <= my_rom(9582); 
 data9 <= my_rom(10937); 
 data10 <= my_rom(12292);
when "00001100010" => 
 data1 <= my_rom(98); 
 data2 <= my_rom(1453); 
 data3 <= my_rom(2808); 
 data4 <= my_rom(4163); 
 data5 <= my_rom(5518); 
 data6 <= my_rom(6873); 
 data7 <= my_rom(8228); 
 data8 <= my_rom(9583); 
 data9 <= my_rom(10938); 
 data10 <= my_rom(12293);
when "00001100011" => 
 data1 <= my_rom(99); 
 data2 <= my_rom(1454); 
 data3 <= my_rom(2809); 
 data4 <= my_rom(4164); 
 data5 <= my_rom(5519); 
 data6 <= my_rom(6874); 
 data7 <= my_rom(8229); 
 data8 <= my_rom(9584); 
 data9 <= my_rom(10939); 
 data10 <= my_rom(12294);
when "00001100100" => 
 data1 <= my_rom(100); 
 data2 <= my_rom(1455); 
 data3 <= my_rom(2810); 
 data4 <= my_rom(4165); 
 data5 <= my_rom(5520); 
 data6 <= my_rom(6875); 
 data7 <= my_rom(8230); 
 data8 <= my_rom(9585); 
 data9 <= my_rom(10940); 
 data10 <= my_rom(12295);
when "00001100101" => 
 data1 <= my_rom(101); 
 data2 <= my_rom(1456); 
 data3 <= my_rom(2811); 
 data4 <= my_rom(4166); 
 data5 <= my_rom(5521); 
 data6 <= my_rom(6876); 
 data7 <= my_rom(8231); 
 data8 <= my_rom(9586); 
 data9 <= my_rom(10941); 
 data10 <= my_rom(12296);
when "00001100110" => 
 data1 <= my_rom(102); 
 data2 <= my_rom(1457); 
 data3 <= my_rom(2812); 
 data4 <= my_rom(4167); 
 data5 <= my_rom(5522); 
 data6 <= my_rom(6877); 
 data7 <= my_rom(8232); 
 data8 <= my_rom(9587); 
 data9 <= my_rom(10942); 
 data10 <= my_rom(12297);
when "00001100111" => 
 data1 <= my_rom(103); 
 data2 <= my_rom(1458); 
 data3 <= my_rom(2813); 
 data4 <= my_rom(4168); 
 data5 <= my_rom(5523); 
 data6 <= my_rom(6878); 
 data7 <= my_rom(8233); 
 data8 <= my_rom(9588); 
 data9 <= my_rom(10943); 
 data10 <= my_rom(12298);
when "00001101000" => 
 data1 <= my_rom(104); 
 data2 <= my_rom(1459); 
 data3 <= my_rom(2814); 
 data4 <= my_rom(4169); 
 data5 <= my_rom(5524); 
 data6 <= my_rom(6879); 
 data7 <= my_rom(8234); 
 data8 <= my_rom(9589); 
 data9 <= my_rom(10944); 
 data10 <= my_rom(12299);
when "00001101001" => 
 data1 <= my_rom(105); 
 data2 <= my_rom(1460); 
 data3 <= my_rom(2815); 
 data4 <= my_rom(4170); 
 data5 <= my_rom(5525); 
 data6 <= my_rom(6880); 
 data7 <= my_rom(8235); 
 data8 <= my_rom(9590); 
 data9 <= my_rom(10945); 
 data10 <= my_rom(12300);
when "00001101010" => 
 data1 <= my_rom(106); 
 data2 <= my_rom(1461); 
 data3 <= my_rom(2816); 
 data4 <= my_rom(4171); 
 data5 <= my_rom(5526); 
 data6 <= my_rom(6881); 
 data7 <= my_rom(8236); 
 data8 <= my_rom(9591); 
 data9 <= my_rom(10946); 
 data10 <= my_rom(12301);
when "00001101011" => 
 data1 <= my_rom(107); 
 data2 <= my_rom(1462); 
 data3 <= my_rom(2817); 
 data4 <= my_rom(4172); 
 data5 <= my_rom(5527); 
 data6 <= my_rom(6882); 
 data7 <= my_rom(8237); 
 data8 <= my_rom(9592); 
 data9 <= my_rom(10947); 
 data10 <= my_rom(12302);
when "00001101100" => 
 data1 <= my_rom(108); 
 data2 <= my_rom(1463); 
 data3 <= my_rom(2818); 
 data4 <= my_rom(4173); 
 data5 <= my_rom(5528); 
 data6 <= my_rom(6883); 
 data7 <= my_rom(8238); 
 data8 <= my_rom(9593); 
 data9 <= my_rom(10948); 
 data10 <= my_rom(12303);
when "00001101101" => 
 data1 <= my_rom(109); 
 data2 <= my_rom(1464); 
 data3 <= my_rom(2819); 
 data4 <= my_rom(4174); 
 data5 <= my_rom(5529); 
 data6 <= my_rom(6884); 
 data7 <= my_rom(8239); 
 data8 <= my_rom(9594); 
 data9 <= my_rom(10949); 
 data10 <= my_rom(12304);
when "00001101110" => 
 data1 <= my_rom(110); 
 data2 <= my_rom(1465); 
 data3 <= my_rom(2820); 
 data4 <= my_rom(4175); 
 data5 <= my_rom(5530); 
 data6 <= my_rom(6885); 
 data7 <= my_rom(8240); 
 data8 <= my_rom(9595); 
 data9 <= my_rom(10950); 
 data10 <= my_rom(12305);
when "00001101111" => 
 data1 <= my_rom(111); 
 data2 <= my_rom(1466); 
 data3 <= my_rom(2821); 
 data4 <= my_rom(4176); 
 data5 <= my_rom(5531); 
 data6 <= my_rom(6886); 
 data7 <= my_rom(8241); 
 data8 <= my_rom(9596); 
 data9 <= my_rom(10951); 
 data10 <= my_rom(12306);
when "00001110000" => 
 data1 <= my_rom(112); 
 data2 <= my_rom(1467); 
 data3 <= my_rom(2822); 
 data4 <= my_rom(4177); 
 data5 <= my_rom(5532); 
 data6 <= my_rom(6887); 
 data7 <= my_rom(8242); 
 data8 <= my_rom(9597); 
 data9 <= my_rom(10952); 
 data10 <= my_rom(12307);
when "00001110001" => 
 data1 <= my_rom(113); 
 data2 <= my_rom(1468); 
 data3 <= my_rom(2823); 
 data4 <= my_rom(4178); 
 data5 <= my_rom(5533); 
 data6 <= my_rom(6888); 
 data7 <= my_rom(8243); 
 data8 <= my_rom(9598); 
 data9 <= my_rom(10953); 
 data10 <= my_rom(12308);
when "00001110010" => 
 data1 <= my_rom(114); 
 data2 <= my_rom(1469); 
 data3 <= my_rom(2824); 
 data4 <= my_rom(4179); 
 data5 <= my_rom(5534); 
 data6 <= my_rom(6889); 
 data7 <= my_rom(8244); 
 data8 <= my_rom(9599); 
 data9 <= my_rom(10954); 
 data10 <= my_rom(12309);
when "00001110011" => 
 data1 <= my_rom(115); 
 data2 <= my_rom(1470); 
 data3 <= my_rom(2825); 
 data4 <= my_rom(4180); 
 data5 <= my_rom(5535); 
 data6 <= my_rom(6890); 
 data7 <= my_rom(8245); 
 data8 <= my_rom(9600); 
 data9 <= my_rom(10955); 
 data10 <= my_rom(12310);
when "00001110100" => 
 data1 <= my_rom(116); 
 data2 <= my_rom(1471); 
 data3 <= my_rom(2826); 
 data4 <= my_rom(4181); 
 data5 <= my_rom(5536); 
 data6 <= my_rom(6891); 
 data7 <= my_rom(8246); 
 data8 <= my_rom(9601); 
 data9 <= my_rom(10956); 
 data10 <= my_rom(12311);
when "00001110101" => 
 data1 <= my_rom(117); 
 data2 <= my_rom(1472); 
 data3 <= my_rom(2827); 
 data4 <= my_rom(4182); 
 data5 <= my_rom(5537); 
 data6 <= my_rom(6892); 
 data7 <= my_rom(8247); 
 data8 <= my_rom(9602); 
 data9 <= my_rom(10957); 
 data10 <= my_rom(12312);
when "00001110110" => 
 data1 <= my_rom(118); 
 data2 <= my_rom(1473); 
 data3 <= my_rom(2828); 
 data4 <= my_rom(4183); 
 data5 <= my_rom(5538); 
 data6 <= my_rom(6893); 
 data7 <= my_rom(8248); 
 data8 <= my_rom(9603); 
 data9 <= my_rom(10958); 
 data10 <= my_rom(12313);
when "00001110111" => 
 data1 <= my_rom(119); 
 data2 <= my_rom(1474); 
 data3 <= my_rom(2829); 
 data4 <= my_rom(4184); 
 data5 <= my_rom(5539); 
 data6 <= my_rom(6894); 
 data7 <= my_rom(8249); 
 data8 <= my_rom(9604); 
 data9 <= my_rom(10959); 
 data10 <= my_rom(12314);
when "00001111000" => 
 data1 <= my_rom(120); 
 data2 <= my_rom(1475); 
 data3 <= my_rom(2830); 
 data4 <= my_rom(4185); 
 data5 <= my_rom(5540); 
 data6 <= my_rom(6895); 
 data7 <= my_rom(8250); 
 data8 <= my_rom(9605); 
 data9 <= my_rom(10960); 
 data10 <= my_rom(12315);
when "00001111001" => 
 data1 <= my_rom(121); 
 data2 <= my_rom(1476); 
 data3 <= my_rom(2831); 
 data4 <= my_rom(4186); 
 data5 <= my_rom(5541); 
 data6 <= my_rom(6896); 
 data7 <= my_rom(8251); 
 data8 <= my_rom(9606); 
 data9 <= my_rom(10961); 
 data10 <= my_rom(12316);
when "00001111010" => 
 data1 <= my_rom(122); 
 data2 <= my_rom(1477); 
 data3 <= my_rom(2832); 
 data4 <= my_rom(4187); 
 data5 <= my_rom(5542); 
 data6 <= my_rom(6897); 
 data7 <= my_rom(8252); 
 data8 <= my_rom(9607); 
 data9 <= my_rom(10962); 
 data10 <= my_rom(12317);
when "00001111011" => 
 data1 <= my_rom(123); 
 data2 <= my_rom(1478); 
 data3 <= my_rom(2833); 
 data4 <= my_rom(4188); 
 data5 <= my_rom(5543); 
 data6 <= my_rom(6898); 
 data7 <= my_rom(8253); 
 data8 <= my_rom(9608); 
 data9 <= my_rom(10963); 
 data10 <= my_rom(12318);
when "00001111100" => 
 data1 <= my_rom(124); 
 data2 <= my_rom(1479); 
 data3 <= my_rom(2834); 
 data4 <= my_rom(4189); 
 data5 <= my_rom(5544); 
 data6 <= my_rom(6899); 
 data7 <= my_rom(8254); 
 data8 <= my_rom(9609); 
 data9 <= my_rom(10964); 
 data10 <= my_rom(12319);
when "00001111101" => 
 data1 <= my_rom(125); 
 data2 <= my_rom(1480); 
 data3 <= my_rom(2835); 
 data4 <= my_rom(4190); 
 data5 <= my_rom(5545); 
 data6 <= my_rom(6900); 
 data7 <= my_rom(8255); 
 data8 <= my_rom(9610); 
 data9 <= my_rom(10965); 
 data10 <= my_rom(12320);
when "00001111110" => 
 data1 <= my_rom(126); 
 data2 <= my_rom(1481); 
 data3 <= my_rom(2836); 
 data4 <= my_rom(4191); 
 data5 <= my_rom(5546); 
 data6 <= my_rom(6901); 
 data7 <= my_rom(8256); 
 data8 <= my_rom(9611); 
 data9 <= my_rom(10966); 
 data10 <= my_rom(12321);
when "00001111111" => 
 data1 <= my_rom(127); 
 data2 <= my_rom(1482); 
 data3 <= my_rom(2837); 
 data4 <= my_rom(4192); 
 data5 <= my_rom(5547); 
 data6 <= my_rom(6902); 
 data7 <= my_rom(8257); 
 data8 <= my_rom(9612); 
 data9 <= my_rom(10967); 
 data10 <= my_rom(12322);
when "00010000000" => 
 data1 <= my_rom(128); 
 data2 <= my_rom(1483); 
 data3 <= my_rom(2838); 
 data4 <= my_rom(4193); 
 data5 <= my_rom(5548); 
 data6 <= my_rom(6903); 
 data7 <= my_rom(8258); 
 data8 <= my_rom(9613); 
 data9 <= my_rom(10968); 
 data10 <= my_rom(12323);
when "00010000001" => 
 data1 <= my_rom(129); 
 data2 <= my_rom(1484); 
 data3 <= my_rom(2839); 
 data4 <= my_rom(4194); 
 data5 <= my_rom(5549); 
 data6 <= my_rom(6904); 
 data7 <= my_rom(8259); 
 data8 <= my_rom(9614); 
 data9 <= my_rom(10969); 
 data10 <= my_rom(12324);
when "00010000010" => 
 data1 <= my_rom(130); 
 data2 <= my_rom(1485); 
 data3 <= my_rom(2840); 
 data4 <= my_rom(4195); 
 data5 <= my_rom(5550); 
 data6 <= my_rom(6905); 
 data7 <= my_rom(8260); 
 data8 <= my_rom(9615); 
 data9 <= my_rom(10970); 
 data10 <= my_rom(12325);
when "00010000011" => 
 data1 <= my_rom(131); 
 data2 <= my_rom(1486); 
 data3 <= my_rom(2841); 
 data4 <= my_rom(4196); 
 data5 <= my_rom(5551); 
 data6 <= my_rom(6906); 
 data7 <= my_rom(8261); 
 data8 <= my_rom(9616); 
 data9 <= my_rom(10971); 
 data10 <= my_rom(12326);
when "00010000100" => 
 data1 <= my_rom(132); 
 data2 <= my_rom(1487); 
 data3 <= my_rom(2842); 
 data4 <= my_rom(4197); 
 data5 <= my_rom(5552); 
 data6 <= my_rom(6907); 
 data7 <= my_rom(8262); 
 data8 <= my_rom(9617); 
 data9 <= my_rom(10972); 
 data10 <= my_rom(12327);
when "00010000101" => 
 data1 <= my_rom(133); 
 data2 <= my_rom(1488); 
 data3 <= my_rom(2843); 
 data4 <= my_rom(4198); 
 data5 <= my_rom(5553); 
 data6 <= my_rom(6908); 
 data7 <= my_rom(8263); 
 data8 <= my_rom(9618); 
 data9 <= my_rom(10973); 
 data10 <= my_rom(12328);
when "00010000110" => 
 data1 <= my_rom(134); 
 data2 <= my_rom(1489); 
 data3 <= my_rom(2844); 
 data4 <= my_rom(4199); 
 data5 <= my_rom(5554); 
 data6 <= my_rom(6909); 
 data7 <= my_rom(8264); 
 data8 <= my_rom(9619); 
 data9 <= my_rom(10974); 
 data10 <= my_rom(12329);
when "00010000111" => 
 data1 <= my_rom(135); 
 data2 <= my_rom(1490); 
 data3 <= my_rom(2845); 
 data4 <= my_rom(4200); 
 data5 <= my_rom(5555); 
 data6 <= my_rom(6910); 
 data7 <= my_rom(8265); 
 data8 <= my_rom(9620); 
 data9 <= my_rom(10975); 
 data10 <= my_rom(12330);
when "00010001000" => 
 data1 <= my_rom(136); 
 data2 <= my_rom(1491); 
 data3 <= my_rom(2846); 
 data4 <= my_rom(4201); 
 data5 <= my_rom(5556); 
 data6 <= my_rom(6911); 
 data7 <= my_rom(8266); 
 data8 <= my_rom(9621); 
 data9 <= my_rom(10976); 
 data10 <= my_rom(12331);
when "00010001001" => 
 data1 <= my_rom(137); 
 data2 <= my_rom(1492); 
 data3 <= my_rom(2847); 
 data4 <= my_rom(4202); 
 data5 <= my_rom(5557); 
 data6 <= my_rom(6912); 
 data7 <= my_rom(8267); 
 data8 <= my_rom(9622); 
 data9 <= my_rom(10977); 
 data10 <= my_rom(12332);
when "00010001010" => 
 data1 <= my_rom(138); 
 data2 <= my_rom(1493); 
 data3 <= my_rom(2848); 
 data4 <= my_rom(4203); 
 data5 <= my_rom(5558); 
 data6 <= my_rom(6913); 
 data7 <= my_rom(8268); 
 data8 <= my_rom(9623); 
 data9 <= my_rom(10978); 
 data10 <= my_rom(12333);
when "00010001011" => 
 data1 <= my_rom(139); 
 data2 <= my_rom(1494); 
 data3 <= my_rom(2849); 
 data4 <= my_rom(4204); 
 data5 <= my_rom(5559); 
 data6 <= my_rom(6914); 
 data7 <= my_rom(8269); 
 data8 <= my_rom(9624); 
 data9 <= my_rom(10979); 
 data10 <= my_rom(12334);
when "00010001100" => 
 data1 <= my_rom(140); 
 data2 <= my_rom(1495); 
 data3 <= my_rom(2850); 
 data4 <= my_rom(4205); 
 data5 <= my_rom(5560); 
 data6 <= my_rom(6915); 
 data7 <= my_rom(8270); 
 data8 <= my_rom(9625); 
 data9 <= my_rom(10980); 
 data10 <= my_rom(12335);
when "00010001101" => 
 data1 <= my_rom(141); 
 data2 <= my_rom(1496); 
 data3 <= my_rom(2851); 
 data4 <= my_rom(4206); 
 data5 <= my_rom(5561); 
 data6 <= my_rom(6916); 
 data7 <= my_rom(8271); 
 data8 <= my_rom(9626); 
 data9 <= my_rom(10981); 
 data10 <= my_rom(12336);
when "00010001110" => 
 data1 <= my_rom(142); 
 data2 <= my_rom(1497); 
 data3 <= my_rom(2852); 
 data4 <= my_rom(4207); 
 data5 <= my_rom(5562); 
 data6 <= my_rom(6917); 
 data7 <= my_rom(8272); 
 data8 <= my_rom(9627); 
 data9 <= my_rom(10982); 
 data10 <= my_rom(12337);
when "00010001111" => 
 data1 <= my_rom(143); 
 data2 <= my_rom(1498); 
 data3 <= my_rom(2853); 
 data4 <= my_rom(4208); 
 data5 <= my_rom(5563); 
 data6 <= my_rom(6918); 
 data7 <= my_rom(8273); 
 data8 <= my_rom(9628); 
 data9 <= my_rom(10983); 
 data10 <= my_rom(12338);
when "00010010000" => 
 data1 <= my_rom(144); 
 data2 <= my_rom(1499); 
 data3 <= my_rom(2854); 
 data4 <= my_rom(4209); 
 data5 <= my_rom(5564); 
 data6 <= my_rom(6919); 
 data7 <= my_rom(8274); 
 data8 <= my_rom(9629); 
 data9 <= my_rom(10984); 
 data10 <= my_rom(12339);
when "00010010001" => 
 data1 <= my_rom(145); 
 data2 <= my_rom(1500); 
 data3 <= my_rom(2855); 
 data4 <= my_rom(4210); 
 data5 <= my_rom(5565); 
 data6 <= my_rom(6920); 
 data7 <= my_rom(8275); 
 data8 <= my_rom(9630); 
 data9 <= my_rom(10985); 
 data10 <= my_rom(12340);
when "00010010010" => 
 data1 <= my_rom(146); 
 data2 <= my_rom(1501); 
 data3 <= my_rom(2856); 
 data4 <= my_rom(4211); 
 data5 <= my_rom(5566); 
 data6 <= my_rom(6921); 
 data7 <= my_rom(8276); 
 data8 <= my_rom(9631); 
 data9 <= my_rom(10986); 
 data10 <= my_rom(12341);
when "00010010011" => 
 data1 <= my_rom(147); 
 data2 <= my_rom(1502); 
 data3 <= my_rom(2857); 
 data4 <= my_rom(4212); 
 data5 <= my_rom(5567); 
 data6 <= my_rom(6922); 
 data7 <= my_rom(8277); 
 data8 <= my_rom(9632); 
 data9 <= my_rom(10987); 
 data10 <= my_rom(12342);
when "00010010100" => 
 data1 <= my_rom(148); 
 data2 <= my_rom(1503); 
 data3 <= my_rom(2858); 
 data4 <= my_rom(4213); 
 data5 <= my_rom(5568); 
 data6 <= my_rom(6923); 
 data7 <= my_rom(8278); 
 data8 <= my_rom(9633); 
 data9 <= my_rom(10988); 
 data10 <= my_rom(12343);
when "00010010101" => 
 data1 <= my_rom(149); 
 data2 <= my_rom(1504); 
 data3 <= my_rom(2859); 
 data4 <= my_rom(4214); 
 data5 <= my_rom(5569); 
 data6 <= my_rom(6924); 
 data7 <= my_rom(8279); 
 data8 <= my_rom(9634); 
 data9 <= my_rom(10989); 
 data10 <= my_rom(12344);
when "00010010110" => 
 data1 <= my_rom(150); 
 data2 <= my_rom(1505); 
 data3 <= my_rom(2860); 
 data4 <= my_rom(4215); 
 data5 <= my_rom(5570); 
 data6 <= my_rom(6925); 
 data7 <= my_rom(8280); 
 data8 <= my_rom(9635); 
 data9 <= my_rom(10990); 
 data10 <= my_rom(12345);
when "00010010111" => 
 data1 <= my_rom(151); 
 data2 <= my_rom(1506); 
 data3 <= my_rom(2861); 
 data4 <= my_rom(4216); 
 data5 <= my_rom(5571); 
 data6 <= my_rom(6926); 
 data7 <= my_rom(8281); 
 data8 <= my_rom(9636); 
 data9 <= my_rom(10991); 
 data10 <= my_rom(12346);
when "00010011000" => 
 data1 <= my_rom(152); 
 data2 <= my_rom(1507); 
 data3 <= my_rom(2862); 
 data4 <= my_rom(4217); 
 data5 <= my_rom(5572); 
 data6 <= my_rom(6927); 
 data7 <= my_rom(8282); 
 data8 <= my_rom(9637); 
 data9 <= my_rom(10992); 
 data10 <= my_rom(12347);
when "00010011001" => 
 data1 <= my_rom(153); 
 data2 <= my_rom(1508); 
 data3 <= my_rom(2863); 
 data4 <= my_rom(4218); 
 data5 <= my_rom(5573); 
 data6 <= my_rom(6928); 
 data7 <= my_rom(8283); 
 data8 <= my_rom(9638); 
 data9 <= my_rom(10993); 
 data10 <= my_rom(12348);
when "00010011010" => 
 data1 <= my_rom(154); 
 data2 <= my_rom(1509); 
 data3 <= my_rom(2864); 
 data4 <= my_rom(4219); 
 data5 <= my_rom(5574); 
 data6 <= my_rom(6929); 
 data7 <= my_rom(8284); 
 data8 <= my_rom(9639); 
 data9 <= my_rom(10994); 
 data10 <= my_rom(12349);
when "00010011011" => 
 data1 <= my_rom(155); 
 data2 <= my_rom(1510); 
 data3 <= my_rom(2865); 
 data4 <= my_rom(4220); 
 data5 <= my_rom(5575); 
 data6 <= my_rom(6930); 
 data7 <= my_rom(8285); 
 data8 <= my_rom(9640); 
 data9 <= my_rom(10995); 
 data10 <= my_rom(12350);
when "00010011100" => 
 data1 <= my_rom(156); 
 data2 <= my_rom(1511); 
 data3 <= my_rom(2866); 
 data4 <= my_rom(4221); 
 data5 <= my_rom(5576); 
 data6 <= my_rom(6931); 
 data7 <= my_rom(8286); 
 data8 <= my_rom(9641); 
 data9 <= my_rom(10996); 
 data10 <= my_rom(12351);
when "00010011101" => 
 data1 <= my_rom(157); 
 data2 <= my_rom(1512); 
 data3 <= my_rom(2867); 
 data4 <= my_rom(4222); 
 data5 <= my_rom(5577); 
 data6 <= my_rom(6932); 
 data7 <= my_rom(8287); 
 data8 <= my_rom(9642); 
 data9 <= my_rom(10997); 
 data10 <= my_rom(12352);
when "00010011110" => 
 data1 <= my_rom(158); 
 data2 <= my_rom(1513); 
 data3 <= my_rom(2868); 
 data4 <= my_rom(4223); 
 data5 <= my_rom(5578); 
 data6 <= my_rom(6933); 
 data7 <= my_rom(8288); 
 data8 <= my_rom(9643); 
 data9 <= my_rom(10998); 
 data10 <= my_rom(12353);
when "00010011111" => 
 data1 <= my_rom(159); 
 data2 <= my_rom(1514); 
 data3 <= my_rom(2869); 
 data4 <= my_rom(4224); 
 data5 <= my_rom(5579); 
 data6 <= my_rom(6934); 
 data7 <= my_rom(8289); 
 data8 <= my_rom(9644); 
 data9 <= my_rom(10999); 
 data10 <= my_rom(12354);
when "00010100000" => 
 data1 <= my_rom(160); 
 data2 <= my_rom(1515); 
 data3 <= my_rom(2870); 
 data4 <= my_rom(4225); 
 data5 <= my_rom(5580); 
 data6 <= my_rom(6935); 
 data7 <= my_rom(8290); 
 data8 <= my_rom(9645); 
 data9 <= my_rom(11000); 
 data10 <= my_rom(12355);
when "00010100001" => 
 data1 <= my_rom(161); 
 data2 <= my_rom(1516); 
 data3 <= my_rom(2871); 
 data4 <= my_rom(4226); 
 data5 <= my_rom(5581); 
 data6 <= my_rom(6936); 
 data7 <= my_rom(8291); 
 data8 <= my_rom(9646); 
 data9 <= my_rom(11001); 
 data10 <= my_rom(12356);
when "00010100010" => 
 data1 <= my_rom(162); 
 data2 <= my_rom(1517); 
 data3 <= my_rom(2872); 
 data4 <= my_rom(4227); 
 data5 <= my_rom(5582); 
 data6 <= my_rom(6937); 
 data7 <= my_rom(8292); 
 data8 <= my_rom(9647); 
 data9 <= my_rom(11002); 
 data10 <= my_rom(12357);
when "00010100011" => 
 data1 <= my_rom(163); 
 data2 <= my_rom(1518); 
 data3 <= my_rom(2873); 
 data4 <= my_rom(4228); 
 data5 <= my_rom(5583); 
 data6 <= my_rom(6938); 
 data7 <= my_rom(8293); 
 data8 <= my_rom(9648); 
 data9 <= my_rom(11003); 
 data10 <= my_rom(12358);
when "00010100100" => 
 data1 <= my_rom(164); 
 data2 <= my_rom(1519); 
 data3 <= my_rom(2874); 
 data4 <= my_rom(4229); 
 data5 <= my_rom(5584); 
 data6 <= my_rom(6939); 
 data7 <= my_rom(8294); 
 data8 <= my_rom(9649); 
 data9 <= my_rom(11004); 
 data10 <= my_rom(12359);
when "00010100101" => 
 data1 <= my_rom(165); 
 data2 <= my_rom(1520); 
 data3 <= my_rom(2875); 
 data4 <= my_rom(4230); 
 data5 <= my_rom(5585); 
 data6 <= my_rom(6940); 
 data7 <= my_rom(8295); 
 data8 <= my_rom(9650); 
 data9 <= my_rom(11005); 
 data10 <= my_rom(12360);
when "00010100110" => 
 data1 <= my_rom(166); 
 data2 <= my_rom(1521); 
 data3 <= my_rom(2876); 
 data4 <= my_rom(4231); 
 data5 <= my_rom(5586); 
 data6 <= my_rom(6941); 
 data7 <= my_rom(8296); 
 data8 <= my_rom(9651); 
 data9 <= my_rom(11006); 
 data10 <= my_rom(12361);
when "00010100111" => 
 data1 <= my_rom(167); 
 data2 <= my_rom(1522); 
 data3 <= my_rom(2877); 
 data4 <= my_rom(4232); 
 data5 <= my_rom(5587); 
 data6 <= my_rom(6942); 
 data7 <= my_rom(8297); 
 data8 <= my_rom(9652); 
 data9 <= my_rom(11007); 
 data10 <= my_rom(12362);
when "00010101000" => 
 data1 <= my_rom(168); 
 data2 <= my_rom(1523); 
 data3 <= my_rom(2878); 
 data4 <= my_rom(4233); 
 data5 <= my_rom(5588); 
 data6 <= my_rom(6943); 
 data7 <= my_rom(8298); 
 data8 <= my_rom(9653); 
 data9 <= my_rom(11008); 
 data10 <= my_rom(12363);
when "00010101001" => 
 data1 <= my_rom(169); 
 data2 <= my_rom(1524); 
 data3 <= my_rom(2879); 
 data4 <= my_rom(4234); 
 data5 <= my_rom(5589); 
 data6 <= my_rom(6944); 
 data7 <= my_rom(8299); 
 data8 <= my_rom(9654); 
 data9 <= my_rom(11009); 
 data10 <= my_rom(12364);
when "00010101010" => 
 data1 <= my_rom(170); 
 data2 <= my_rom(1525); 
 data3 <= my_rom(2880); 
 data4 <= my_rom(4235); 
 data5 <= my_rom(5590); 
 data6 <= my_rom(6945); 
 data7 <= my_rom(8300); 
 data8 <= my_rom(9655); 
 data9 <= my_rom(11010); 
 data10 <= my_rom(12365);
when "00010101011" => 
 data1 <= my_rom(171); 
 data2 <= my_rom(1526); 
 data3 <= my_rom(2881); 
 data4 <= my_rom(4236); 
 data5 <= my_rom(5591); 
 data6 <= my_rom(6946); 
 data7 <= my_rom(8301); 
 data8 <= my_rom(9656); 
 data9 <= my_rom(11011); 
 data10 <= my_rom(12366);
when "00010101100" => 
 data1 <= my_rom(172); 
 data2 <= my_rom(1527); 
 data3 <= my_rom(2882); 
 data4 <= my_rom(4237); 
 data5 <= my_rom(5592); 
 data6 <= my_rom(6947); 
 data7 <= my_rom(8302); 
 data8 <= my_rom(9657); 
 data9 <= my_rom(11012); 
 data10 <= my_rom(12367);
when "00010101101" => 
 data1 <= my_rom(173); 
 data2 <= my_rom(1528); 
 data3 <= my_rom(2883); 
 data4 <= my_rom(4238); 
 data5 <= my_rom(5593); 
 data6 <= my_rom(6948); 
 data7 <= my_rom(8303); 
 data8 <= my_rom(9658); 
 data9 <= my_rom(11013); 
 data10 <= my_rom(12368);
when "00010101110" => 
 data1 <= my_rom(174); 
 data2 <= my_rom(1529); 
 data3 <= my_rom(2884); 
 data4 <= my_rom(4239); 
 data5 <= my_rom(5594); 
 data6 <= my_rom(6949); 
 data7 <= my_rom(8304); 
 data8 <= my_rom(9659); 
 data9 <= my_rom(11014); 
 data10 <= my_rom(12369);
when "00010101111" => 
 data1 <= my_rom(175); 
 data2 <= my_rom(1530); 
 data3 <= my_rom(2885); 
 data4 <= my_rom(4240); 
 data5 <= my_rom(5595); 
 data6 <= my_rom(6950); 
 data7 <= my_rom(8305); 
 data8 <= my_rom(9660); 
 data9 <= my_rom(11015); 
 data10 <= my_rom(12370);
when "00010110000" => 
 data1 <= my_rom(176); 
 data2 <= my_rom(1531); 
 data3 <= my_rom(2886); 
 data4 <= my_rom(4241); 
 data5 <= my_rom(5596); 
 data6 <= my_rom(6951); 
 data7 <= my_rom(8306); 
 data8 <= my_rom(9661); 
 data9 <= my_rom(11016); 
 data10 <= my_rom(12371);
when "00010110001" => 
 data1 <= my_rom(177); 
 data2 <= my_rom(1532); 
 data3 <= my_rom(2887); 
 data4 <= my_rom(4242); 
 data5 <= my_rom(5597); 
 data6 <= my_rom(6952); 
 data7 <= my_rom(8307); 
 data8 <= my_rom(9662); 
 data9 <= my_rom(11017); 
 data10 <= my_rom(12372);
when "00010110010" => 
 data1 <= my_rom(178); 
 data2 <= my_rom(1533); 
 data3 <= my_rom(2888); 
 data4 <= my_rom(4243); 
 data5 <= my_rom(5598); 
 data6 <= my_rom(6953); 
 data7 <= my_rom(8308); 
 data8 <= my_rom(9663); 
 data9 <= my_rom(11018); 
 data10 <= my_rom(12373);
when "00010110011" => 
 data1 <= my_rom(179); 
 data2 <= my_rom(1534); 
 data3 <= my_rom(2889); 
 data4 <= my_rom(4244); 
 data5 <= my_rom(5599); 
 data6 <= my_rom(6954); 
 data7 <= my_rom(8309); 
 data8 <= my_rom(9664); 
 data9 <= my_rom(11019); 
 data10 <= my_rom(12374);
when "00010110100" => 
 data1 <= my_rom(180); 
 data2 <= my_rom(1535); 
 data3 <= my_rom(2890); 
 data4 <= my_rom(4245); 
 data5 <= my_rom(5600); 
 data6 <= my_rom(6955); 
 data7 <= my_rom(8310); 
 data8 <= my_rom(9665); 
 data9 <= my_rom(11020); 
 data10 <= my_rom(12375);
when "00010110101" => 
 data1 <= my_rom(181); 
 data2 <= my_rom(1536); 
 data3 <= my_rom(2891); 
 data4 <= my_rom(4246); 
 data5 <= my_rom(5601); 
 data6 <= my_rom(6956); 
 data7 <= my_rom(8311); 
 data8 <= my_rom(9666); 
 data9 <= my_rom(11021); 
 data10 <= my_rom(12376);
when "00010110110" => 
 data1 <= my_rom(182); 
 data2 <= my_rom(1537); 
 data3 <= my_rom(2892); 
 data4 <= my_rom(4247); 
 data5 <= my_rom(5602); 
 data6 <= my_rom(6957); 
 data7 <= my_rom(8312); 
 data8 <= my_rom(9667); 
 data9 <= my_rom(11022); 
 data10 <= my_rom(12377);
when "00010110111" => 
 data1 <= my_rom(183); 
 data2 <= my_rom(1538); 
 data3 <= my_rom(2893); 
 data4 <= my_rom(4248); 
 data5 <= my_rom(5603); 
 data6 <= my_rom(6958); 
 data7 <= my_rom(8313); 
 data8 <= my_rom(9668); 
 data9 <= my_rom(11023); 
 data10 <= my_rom(12378);
when "00010111000" => 
 data1 <= my_rom(184); 
 data2 <= my_rom(1539); 
 data3 <= my_rom(2894); 
 data4 <= my_rom(4249); 
 data5 <= my_rom(5604); 
 data6 <= my_rom(6959); 
 data7 <= my_rom(8314); 
 data8 <= my_rom(9669); 
 data9 <= my_rom(11024); 
 data10 <= my_rom(12379);
when "00010111001" => 
 data1 <= my_rom(185); 
 data2 <= my_rom(1540); 
 data3 <= my_rom(2895); 
 data4 <= my_rom(4250); 
 data5 <= my_rom(5605); 
 data6 <= my_rom(6960); 
 data7 <= my_rom(8315); 
 data8 <= my_rom(9670); 
 data9 <= my_rom(11025); 
 data10 <= my_rom(12380);
when "00010111010" => 
 data1 <= my_rom(186); 
 data2 <= my_rom(1541); 
 data3 <= my_rom(2896); 
 data4 <= my_rom(4251); 
 data5 <= my_rom(5606); 
 data6 <= my_rom(6961); 
 data7 <= my_rom(8316); 
 data8 <= my_rom(9671); 
 data9 <= my_rom(11026); 
 data10 <= my_rom(12381);
when "00010111011" => 
 data1 <= my_rom(187); 
 data2 <= my_rom(1542); 
 data3 <= my_rom(2897); 
 data4 <= my_rom(4252); 
 data5 <= my_rom(5607); 
 data6 <= my_rom(6962); 
 data7 <= my_rom(8317); 
 data8 <= my_rom(9672); 
 data9 <= my_rom(11027); 
 data10 <= my_rom(12382);
when "00010111100" => 
 data1 <= my_rom(188); 
 data2 <= my_rom(1543); 
 data3 <= my_rom(2898); 
 data4 <= my_rom(4253); 
 data5 <= my_rom(5608); 
 data6 <= my_rom(6963); 
 data7 <= my_rom(8318); 
 data8 <= my_rom(9673); 
 data9 <= my_rom(11028); 
 data10 <= my_rom(12383);
when "00010111101" => 
 data1 <= my_rom(189); 
 data2 <= my_rom(1544); 
 data3 <= my_rom(2899); 
 data4 <= my_rom(4254); 
 data5 <= my_rom(5609); 
 data6 <= my_rom(6964); 
 data7 <= my_rom(8319); 
 data8 <= my_rom(9674); 
 data9 <= my_rom(11029); 
 data10 <= my_rom(12384);
when "00010111110" => 
 data1 <= my_rom(190); 
 data2 <= my_rom(1545); 
 data3 <= my_rom(2900); 
 data4 <= my_rom(4255); 
 data5 <= my_rom(5610); 
 data6 <= my_rom(6965); 
 data7 <= my_rom(8320); 
 data8 <= my_rom(9675); 
 data9 <= my_rom(11030); 
 data10 <= my_rom(12385);
when "00010111111" => 
 data1 <= my_rom(191); 
 data2 <= my_rom(1546); 
 data3 <= my_rom(2901); 
 data4 <= my_rom(4256); 
 data5 <= my_rom(5611); 
 data6 <= my_rom(6966); 
 data7 <= my_rom(8321); 
 data8 <= my_rom(9676); 
 data9 <= my_rom(11031); 
 data10 <= my_rom(12386);
when "00011000000" => 
 data1 <= my_rom(192); 
 data2 <= my_rom(1547); 
 data3 <= my_rom(2902); 
 data4 <= my_rom(4257); 
 data5 <= my_rom(5612); 
 data6 <= my_rom(6967); 
 data7 <= my_rom(8322); 
 data8 <= my_rom(9677); 
 data9 <= my_rom(11032); 
 data10 <= my_rom(12387);
when "00011000001" => 
 data1 <= my_rom(193); 
 data2 <= my_rom(1548); 
 data3 <= my_rom(2903); 
 data4 <= my_rom(4258); 
 data5 <= my_rom(5613); 
 data6 <= my_rom(6968); 
 data7 <= my_rom(8323); 
 data8 <= my_rom(9678); 
 data9 <= my_rom(11033); 
 data10 <= my_rom(12388);
when "00011000010" => 
 data1 <= my_rom(194); 
 data2 <= my_rom(1549); 
 data3 <= my_rom(2904); 
 data4 <= my_rom(4259); 
 data5 <= my_rom(5614); 
 data6 <= my_rom(6969); 
 data7 <= my_rom(8324); 
 data8 <= my_rom(9679); 
 data9 <= my_rom(11034); 
 data10 <= my_rom(12389);
when "00011000011" => 
 data1 <= my_rom(195); 
 data2 <= my_rom(1550); 
 data3 <= my_rom(2905); 
 data4 <= my_rom(4260); 
 data5 <= my_rom(5615); 
 data6 <= my_rom(6970); 
 data7 <= my_rom(8325); 
 data8 <= my_rom(9680); 
 data9 <= my_rom(11035); 
 data10 <= my_rom(12390);
when "00011000100" => 
 data1 <= my_rom(196); 
 data2 <= my_rom(1551); 
 data3 <= my_rom(2906); 
 data4 <= my_rom(4261); 
 data5 <= my_rom(5616); 
 data6 <= my_rom(6971); 
 data7 <= my_rom(8326); 
 data8 <= my_rom(9681); 
 data9 <= my_rom(11036); 
 data10 <= my_rom(12391);
when "00011000101" => 
 data1 <= my_rom(197); 
 data2 <= my_rom(1552); 
 data3 <= my_rom(2907); 
 data4 <= my_rom(4262); 
 data5 <= my_rom(5617); 
 data6 <= my_rom(6972); 
 data7 <= my_rom(8327); 
 data8 <= my_rom(9682); 
 data9 <= my_rom(11037); 
 data10 <= my_rom(12392);
when "00011000110" => 
 data1 <= my_rom(198); 
 data2 <= my_rom(1553); 
 data3 <= my_rom(2908); 
 data4 <= my_rom(4263); 
 data5 <= my_rom(5618); 
 data6 <= my_rom(6973); 
 data7 <= my_rom(8328); 
 data8 <= my_rom(9683); 
 data9 <= my_rom(11038); 
 data10 <= my_rom(12393);
when "00011000111" => 
 data1 <= my_rom(199); 
 data2 <= my_rom(1554); 
 data3 <= my_rom(2909); 
 data4 <= my_rom(4264); 
 data5 <= my_rom(5619); 
 data6 <= my_rom(6974); 
 data7 <= my_rom(8329); 
 data8 <= my_rom(9684); 
 data9 <= my_rom(11039); 
 data10 <= my_rom(12394);
when "00011001000" => 
 data1 <= my_rom(200); 
 data2 <= my_rom(1555); 
 data3 <= my_rom(2910); 
 data4 <= my_rom(4265); 
 data5 <= my_rom(5620); 
 data6 <= my_rom(6975); 
 data7 <= my_rom(8330); 
 data8 <= my_rom(9685); 
 data9 <= my_rom(11040); 
 data10 <= my_rom(12395);
when "00011001001" => 
 data1 <= my_rom(201); 
 data2 <= my_rom(1556); 
 data3 <= my_rom(2911); 
 data4 <= my_rom(4266); 
 data5 <= my_rom(5621); 
 data6 <= my_rom(6976); 
 data7 <= my_rom(8331); 
 data8 <= my_rom(9686); 
 data9 <= my_rom(11041); 
 data10 <= my_rom(12396);
when "00011001010" => 
 data1 <= my_rom(202); 
 data2 <= my_rom(1557); 
 data3 <= my_rom(2912); 
 data4 <= my_rom(4267); 
 data5 <= my_rom(5622); 
 data6 <= my_rom(6977); 
 data7 <= my_rom(8332); 
 data8 <= my_rom(9687); 
 data9 <= my_rom(11042); 
 data10 <= my_rom(12397);
when "00011001011" => 
 data1 <= my_rom(203); 
 data2 <= my_rom(1558); 
 data3 <= my_rom(2913); 
 data4 <= my_rom(4268); 
 data5 <= my_rom(5623); 
 data6 <= my_rom(6978); 
 data7 <= my_rom(8333); 
 data8 <= my_rom(9688); 
 data9 <= my_rom(11043); 
 data10 <= my_rom(12398);
when "00011001100" => 
 data1 <= my_rom(204); 
 data2 <= my_rom(1559); 
 data3 <= my_rom(2914); 
 data4 <= my_rom(4269); 
 data5 <= my_rom(5624); 
 data6 <= my_rom(6979); 
 data7 <= my_rom(8334); 
 data8 <= my_rom(9689); 
 data9 <= my_rom(11044); 
 data10 <= my_rom(12399);
when "00011001101" => 
 data1 <= my_rom(205); 
 data2 <= my_rom(1560); 
 data3 <= my_rom(2915); 
 data4 <= my_rom(4270); 
 data5 <= my_rom(5625); 
 data6 <= my_rom(6980); 
 data7 <= my_rom(8335); 
 data8 <= my_rom(9690); 
 data9 <= my_rom(11045); 
 data10 <= my_rom(12400);
when "00011001110" => 
 data1 <= my_rom(206); 
 data2 <= my_rom(1561); 
 data3 <= my_rom(2916); 
 data4 <= my_rom(4271); 
 data5 <= my_rom(5626); 
 data6 <= my_rom(6981); 
 data7 <= my_rom(8336); 
 data8 <= my_rom(9691); 
 data9 <= my_rom(11046); 
 data10 <= my_rom(12401);
when "00011001111" => 
 data1 <= my_rom(207); 
 data2 <= my_rom(1562); 
 data3 <= my_rom(2917); 
 data4 <= my_rom(4272); 
 data5 <= my_rom(5627); 
 data6 <= my_rom(6982); 
 data7 <= my_rom(8337); 
 data8 <= my_rom(9692); 
 data9 <= my_rom(11047); 
 data10 <= my_rom(12402);
when "00011010000" => 
 data1 <= my_rom(208); 
 data2 <= my_rom(1563); 
 data3 <= my_rom(2918); 
 data4 <= my_rom(4273); 
 data5 <= my_rom(5628); 
 data6 <= my_rom(6983); 
 data7 <= my_rom(8338); 
 data8 <= my_rom(9693); 
 data9 <= my_rom(11048); 
 data10 <= my_rom(12403);
when "00011010001" => 
 data1 <= my_rom(209); 
 data2 <= my_rom(1564); 
 data3 <= my_rom(2919); 
 data4 <= my_rom(4274); 
 data5 <= my_rom(5629); 
 data6 <= my_rom(6984); 
 data7 <= my_rom(8339); 
 data8 <= my_rom(9694); 
 data9 <= my_rom(11049); 
 data10 <= my_rom(12404);
when "00011010010" => 
 data1 <= my_rom(210); 
 data2 <= my_rom(1565); 
 data3 <= my_rom(2920); 
 data4 <= my_rom(4275); 
 data5 <= my_rom(5630); 
 data6 <= my_rom(6985); 
 data7 <= my_rom(8340); 
 data8 <= my_rom(9695); 
 data9 <= my_rom(11050); 
 data10 <= my_rom(12405);
when "00011010011" => 
 data1 <= my_rom(211); 
 data2 <= my_rom(1566); 
 data3 <= my_rom(2921); 
 data4 <= my_rom(4276); 
 data5 <= my_rom(5631); 
 data6 <= my_rom(6986); 
 data7 <= my_rom(8341); 
 data8 <= my_rom(9696); 
 data9 <= my_rom(11051); 
 data10 <= my_rom(12406);
when "00011010100" => 
 data1 <= my_rom(212); 
 data2 <= my_rom(1567); 
 data3 <= my_rom(2922); 
 data4 <= my_rom(4277); 
 data5 <= my_rom(5632); 
 data6 <= my_rom(6987); 
 data7 <= my_rom(8342); 
 data8 <= my_rom(9697); 
 data9 <= my_rom(11052); 
 data10 <= my_rom(12407);
when "00011010101" => 
 data1 <= my_rom(213); 
 data2 <= my_rom(1568); 
 data3 <= my_rom(2923); 
 data4 <= my_rom(4278); 
 data5 <= my_rom(5633); 
 data6 <= my_rom(6988); 
 data7 <= my_rom(8343); 
 data8 <= my_rom(9698); 
 data9 <= my_rom(11053); 
 data10 <= my_rom(12408);
when "00011010110" => 
 data1 <= my_rom(214); 
 data2 <= my_rom(1569); 
 data3 <= my_rom(2924); 
 data4 <= my_rom(4279); 
 data5 <= my_rom(5634); 
 data6 <= my_rom(6989); 
 data7 <= my_rom(8344); 
 data8 <= my_rom(9699); 
 data9 <= my_rom(11054); 
 data10 <= my_rom(12409);
when "00011010111" => 
 data1 <= my_rom(215); 
 data2 <= my_rom(1570); 
 data3 <= my_rom(2925); 
 data4 <= my_rom(4280); 
 data5 <= my_rom(5635); 
 data6 <= my_rom(6990); 
 data7 <= my_rom(8345); 
 data8 <= my_rom(9700); 
 data9 <= my_rom(11055); 
 data10 <= my_rom(12410);
when "00011011000" => 
 data1 <= my_rom(216); 
 data2 <= my_rom(1571); 
 data3 <= my_rom(2926); 
 data4 <= my_rom(4281); 
 data5 <= my_rom(5636); 
 data6 <= my_rom(6991); 
 data7 <= my_rom(8346); 
 data8 <= my_rom(9701); 
 data9 <= my_rom(11056); 
 data10 <= my_rom(12411);
when "00011011001" => 
 data1 <= my_rom(217); 
 data2 <= my_rom(1572); 
 data3 <= my_rom(2927); 
 data4 <= my_rom(4282); 
 data5 <= my_rom(5637); 
 data6 <= my_rom(6992); 
 data7 <= my_rom(8347); 
 data8 <= my_rom(9702); 
 data9 <= my_rom(11057); 
 data10 <= my_rom(12412);
when "00011011010" => 
 data1 <= my_rom(218); 
 data2 <= my_rom(1573); 
 data3 <= my_rom(2928); 
 data4 <= my_rom(4283); 
 data5 <= my_rom(5638); 
 data6 <= my_rom(6993); 
 data7 <= my_rom(8348); 
 data8 <= my_rom(9703); 
 data9 <= my_rom(11058); 
 data10 <= my_rom(12413);
when "00011011011" => 
 data1 <= my_rom(219); 
 data2 <= my_rom(1574); 
 data3 <= my_rom(2929); 
 data4 <= my_rom(4284); 
 data5 <= my_rom(5639); 
 data6 <= my_rom(6994); 
 data7 <= my_rom(8349); 
 data8 <= my_rom(9704); 
 data9 <= my_rom(11059); 
 data10 <= my_rom(12414);
when "00011011100" => 
 data1 <= my_rom(220); 
 data2 <= my_rom(1575); 
 data3 <= my_rom(2930); 
 data4 <= my_rom(4285); 
 data5 <= my_rom(5640); 
 data6 <= my_rom(6995); 
 data7 <= my_rom(8350); 
 data8 <= my_rom(9705); 
 data9 <= my_rom(11060); 
 data10 <= my_rom(12415);
when "00011011101" => 
 data1 <= my_rom(221); 
 data2 <= my_rom(1576); 
 data3 <= my_rom(2931); 
 data4 <= my_rom(4286); 
 data5 <= my_rom(5641); 
 data6 <= my_rom(6996); 
 data7 <= my_rom(8351); 
 data8 <= my_rom(9706); 
 data9 <= my_rom(11061); 
 data10 <= my_rom(12416);
when "00011011110" => 
 data1 <= my_rom(222); 
 data2 <= my_rom(1577); 
 data3 <= my_rom(2932); 
 data4 <= my_rom(4287); 
 data5 <= my_rom(5642); 
 data6 <= my_rom(6997); 
 data7 <= my_rom(8352); 
 data8 <= my_rom(9707); 
 data9 <= my_rom(11062); 
 data10 <= my_rom(12417);
when "00011011111" => 
 data1 <= my_rom(223); 
 data2 <= my_rom(1578); 
 data3 <= my_rom(2933); 
 data4 <= my_rom(4288); 
 data5 <= my_rom(5643); 
 data6 <= my_rom(6998); 
 data7 <= my_rom(8353); 
 data8 <= my_rom(9708); 
 data9 <= my_rom(11063); 
 data10 <= my_rom(12418);
when "00011100000" => 
 data1 <= my_rom(224); 
 data2 <= my_rom(1579); 
 data3 <= my_rom(2934); 
 data4 <= my_rom(4289); 
 data5 <= my_rom(5644); 
 data6 <= my_rom(6999); 
 data7 <= my_rom(8354); 
 data8 <= my_rom(9709); 
 data9 <= my_rom(11064); 
 data10 <= my_rom(12419);
when "00011100001" => 
 data1 <= my_rom(225); 
 data2 <= my_rom(1580); 
 data3 <= my_rom(2935); 
 data4 <= my_rom(4290); 
 data5 <= my_rom(5645); 
 data6 <= my_rom(7000); 
 data7 <= my_rom(8355); 
 data8 <= my_rom(9710); 
 data9 <= my_rom(11065); 
 data10 <= my_rom(12420);
when "00011100010" => 
 data1 <= my_rom(226); 
 data2 <= my_rom(1581); 
 data3 <= my_rom(2936); 
 data4 <= my_rom(4291); 
 data5 <= my_rom(5646); 
 data6 <= my_rom(7001); 
 data7 <= my_rom(8356); 
 data8 <= my_rom(9711); 
 data9 <= my_rom(11066); 
 data10 <= my_rom(12421);
when "00011100011" => 
 data1 <= my_rom(227); 
 data2 <= my_rom(1582); 
 data3 <= my_rom(2937); 
 data4 <= my_rom(4292); 
 data5 <= my_rom(5647); 
 data6 <= my_rom(7002); 
 data7 <= my_rom(8357); 
 data8 <= my_rom(9712); 
 data9 <= my_rom(11067); 
 data10 <= my_rom(12422);
when "00011100100" => 
 data1 <= my_rom(228); 
 data2 <= my_rom(1583); 
 data3 <= my_rom(2938); 
 data4 <= my_rom(4293); 
 data5 <= my_rom(5648); 
 data6 <= my_rom(7003); 
 data7 <= my_rom(8358); 
 data8 <= my_rom(9713); 
 data9 <= my_rom(11068); 
 data10 <= my_rom(12423);
when "00011100101" => 
 data1 <= my_rom(229); 
 data2 <= my_rom(1584); 
 data3 <= my_rom(2939); 
 data4 <= my_rom(4294); 
 data5 <= my_rom(5649); 
 data6 <= my_rom(7004); 
 data7 <= my_rom(8359); 
 data8 <= my_rom(9714); 
 data9 <= my_rom(11069); 
 data10 <= my_rom(12424);
when "00011100110" => 
 data1 <= my_rom(230); 
 data2 <= my_rom(1585); 
 data3 <= my_rom(2940); 
 data4 <= my_rom(4295); 
 data5 <= my_rom(5650); 
 data6 <= my_rom(7005); 
 data7 <= my_rom(8360); 
 data8 <= my_rom(9715); 
 data9 <= my_rom(11070); 
 data10 <= my_rom(12425);
when "00011100111" => 
 data1 <= my_rom(231); 
 data2 <= my_rom(1586); 
 data3 <= my_rom(2941); 
 data4 <= my_rom(4296); 
 data5 <= my_rom(5651); 
 data6 <= my_rom(7006); 
 data7 <= my_rom(8361); 
 data8 <= my_rom(9716); 
 data9 <= my_rom(11071); 
 data10 <= my_rom(12426);
when "00011101000" => 
 data1 <= my_rom(232); 
 data2 <= my_rom(1587); 
 data3 <= my_rom(2942); 
 data4 <= my_rom(4297); 
 data5 <= my_rom(5652); 
 data6 <= my_rom(7007); 
 data7 <= my_rom(8362); 
 data8 <= my_rom(9717); 
 data9 <= my_rom(11072); 
 data10 <= my_rom(12427);
when "00011101001" => 
 data1 <= my_rom(233); 
 data2 <= my_rom(1588); 
 data3 <= my_rom(2943); 
 data4 <= my_rom(4298); 
 data5 <= my_rom(5653); 
 data6 <= my_rom(7008); 
 data7 <= my_rom(8363); 
 data8 <= my_rom(9718); 
 data9 <= my_rom(11073); 
 data10 <= my_rom(12428);
when "00011101010" => 
 data1 <= my_rom(234); 
 data2 <= my_rom(1589); 
 data3 <= my_rom(2944); 
 data4 <= my_rom(4299); 
 data5 <= my_rom(5654); 
 data6 <= my_rom(7009); 
 data7 <= my_rom(8364); 
 data8 <= my_rom(9719); 
 data9 <= my_rom(11074); 
 data10 <= my_rom(12429);
when "00011101011" => 
 data1 <= my_rom(235); 
 data2 <= my_rom(1590); 
 data3 <= my_rom(2945); 
 data4 <= my_rom(4300); 
 data5 <= my_rom(5655); 
 data6 <= my_rom(7010); 
 data7 <= my_rom(8365); 
 data8 <= my_rom(9720); 
 data9 <= my_rom(11075); 
 data10 <= my_rom(12430);
when "00011101100" => 
 data1 <= my_rom(236); 
 data2 <= my_rom(1591); 
 data3 <= my_rom(2946); 
 data4 <= my_rom(4301); 
 data5 <= my_rom(5656); 
 data6 <= my_rom(7011); 
 data7 <= my_rom(8366); 
 data8 <= my_rom(9721); 
 data9 <= my_rom(11076); 
 data10 <= my_rom(12431);
when "00011101101" => 
 data1 <= my_rom(237); 
 data2 <= my_rom(1592); 
 data3 <= my_rom(2947); 
 data4 <= my_rom(4302); 
 data5 <= my_rom(5657); 
 data6 <= my_rom(7012); 
 data7 <= my_rom(8367); 
 data8 <= my_rom(9722); 
 data9 <= my_rom(11077); 
 data10 <= my_rom(12432);
when "00011101110" => 
 data1 <= my_rom(238); 
 data2 <= my_rom(1593); 
 data3 <= my_rom(2948); 
 data4 <= my_rom(4303); 
 data5 <= my_rom(5658); 
 data6 <= my_rom(7013); 
 data7 <= my_rom(8368); 
 data8 <= my_rom(9723); 
 data9 <= my_rom(11078); 
 data10 <= my_rom(12433);
when "00011101111" => 
 data1 <= my_rom(239); 
 data2 <= my_rom(1594); 
 data3 <= my_rom(2949); 
 data4 <= my_rom(4304); 
 data5 <= my_rom(5659); 
 data6 <= my_rom(7014); 
 data7 <= my_rom(8369); 
 data8 <= my_rom(9724); 
 data9 <= my_rom(11079); 
 data10 <= my_rom(12434);
when "00011110000" => 
 data1 <= my_rom(240); 
 data2 <= my_rom(1595); 
 data3 <= my_rom(2950); 
 data4 <= my_rom(4305); 
 data5 <= my_rom(5660); 
 data6 <= my_rom(7015); 
 data7 <= my_rom(8370); 
 data8 <= my_rom(9725); 
 data9 <= my_rom(11080); 
 data10 <= my_rom(12435);
when "00011110001" => 
 data1 <= my_rom(241); 
 data2 <= my_rom(1596); 
 data3 <= my_rom(2951); 
 data4 <= my_rom(4306); 
 data5 <= my_rom(5661); 
 data6 <= my_rom(7016); 
 data7 <= my_rom(8371); 
 data8 <= my_rom(9726); 
 data9 <= my_rom(11081); 
 data10 <= my_rom(12436);
when "00011110010" => 
 data1 <= my_rom(242); 
 data2 <= my_rom(1597); 
 data3 <= my_rom(2952); 
 data4 <= my_rom(4307); 
 data5 <= my_rom(5662); 
 data6 <= my_rom(7017); 
 data7 <= my_rom(8372); 
 data8 <= my_rom(9727); 
 data9 <= my_rom(11082); 
 data10 <= my_rom(12437);
when "00011110011" => 
 data1 <= my_rom(243); 
 data2 <= my_rom(1598); 
 data3 <= my_rom(2953); 
 data4 <= my_rom(4308); 
 data5 <= my_rom(5663); 
 data6 <= my_rom(7018); 
 data7 <= my_rom(8373); 
 data8 <= my_rom(9728); 
 data9 <= my_rom(11083); 
 data10 <= my_rom(12438);
when "00011110100" => 
 data1 <= my_rom(244); 
 data2 <= my_rom(1599); 
 data3 <= my_rom(2954); 
 data4 <= my_rom(4309); 
 data5 <= my_rom(5664); 
 data6 <= my_rom(7019); 
 data7 <= my_rom(8374); 
 data8 <= my_rom(9729); 
 data9 <= my_rom(11084); 
 data10 <= my_rom(12439);
when "00011110101" => 
 data1 <= my_rom(245); 
 data2 <= my_rom(1600); 
 data3 <= my_rom(2955); 
 data4 <= my_rom(4310); 
 data5 <= my_rom(5665); 
 data6 <= my_rom(7020); 
 data7 <= my_rom(8375); 
 data8 <= my_rom(9730); 
 data9 <= my_rom(11085); 
 data10 <= my_rom(12440);
when "00011110110" => 
 data1 <= my_rom(246); 
 data2 <= my_rom(1601); 
 data3 <= my_rom(2956); 
 data4 <= my_rom(4311); 
 data5 <= my_rom(5666); 
 data6 <= my_rom(7021); 
 data7 <= my_rom(8376); 
 data8 <= my_rom(9731); 
 data9 <= my_rom(11086); 
 data10 <= my_rom(12441);
when "00011110111" => 
 data1 <= my_rom(247); 
 data2 <= my_rom(1602); 
 data3 <= my_rom(2957); 
 data4 <= my_rom(4312); 
 data5 <= my_rom(5667); 
 data6 <= my_rom(7022); 
 data7 <= my_rom(8377); 
 data8 <= my_rom(9732); 
 data9 <= my_rom(11087); 
 data10 <= my_rom(12442);
when "00011111000" => 
 data1 <= my_rom(248); 
 data2 <= my_rom(1603); 
 data3 <= my_rom(2958); 
 data4 <= my_rom(4313); 
 data5 <= my_rom(5668); 
 data6 <= my_rom(7023); 
 data7 <= my_rom(8378); 
 data8 <= my_rom(9733); 
 data9 <= my_rom(11088); 
 data10 <= my_rom(12443);
when "00011111001" => 
 data1 <= my_rom(249); 
 data2 <= my_rom(1604); 
 data3 <= my_rom(2959); 
 data4 <= my_rom(4314); 
 data5 <= my_rom(5669); 
 data6 <= my_rom(7024); 
 data7 <= my_rom(8379); 
 data8 <= my_rom(9734); 
 data9 <= my_rom(11089); 
 data10 <= my_rom(12444);
when "00011111010" => 
 data1 <= my_rom(250); 
 data2 <= my_rom(1605); 
 data3 <= my_rom(2960); 
 data4 <= my_rom(4315); 
 data5 <= my_rom(5670); 
 data6 <= my_rom(7025); 
 data7 <= my_rom(8380); 
 data8 <= my_rom(9735); 
 data9 <= my_rom(11090); 
 data10 <= my_rom(12445);
when "00011111011" => 
 data1 <= my_rom(251); 
 data2 <= my_rom(1606); 
 data3 <= my_rom(2961); 
 data4 <= my_rom(4316); 
 data5 <= my_rom(5671); 
 data6 <= my_rom(7026); 
 data7 <= my_rom(8381); 
 data8 <= my_rom(9736); 
 data9 <= my_rom(11091); 
 data10 <= my_rom(12446);
when "00011111100" => 
 data1 <= my_rom(252); 
 data2 <= my_rom(1607); 
 data3 <= my_rom(2962); 
 data4 <= my_rom(4317); 
 data5 <= my_rom(5672); 
 data6 <= my_rom(7027); 
 data7 <= my_rom(8382); 
 data8 <= my_rom(9737); 
 data9 <= my_rom(11092); 
 data10 <= my_rom(12447);
when "00011111101" => 
 data1 <= my_rom(253); 
 data2 <= my_rom(1608); 
 data3 <= my_rom(2963); 
 data4 <= my_rom(4318); 
 data5 <= my_rom(5673); 
 data6 <= my_rom(7028); 
 data7 <= my_rom(8383); 
 data8 <= my_rom(9738); 
 data9 <= my_rom(11093); 
 data10 <= my_rom(12448);
when "00011111110" => 
 data1 <= my_rom(254); 
 data2 <= my_rom(1609); 
 data3 <= my_rom(2964); 
 data4 <= my_rom(4319); 
 data5 <= my_rom(5674); 
 data6 <= my_rom(7029); 
 data7 <= my_rom(8384); 
 data8 <= my_rom(9739); 
 data9 <= my_rom(11094); 
 data10 <= my_rom(12449);
when "00011111111" => 
 data1 <= my_rom(255); 
 data2 <= my_rom(1610); 
 data3 <= my_rom(2965); 
 data4 <= my_rom(4320); 
 data5 <= my_rom(5675); 
 data6 <= my_rom(7030); 
 data7 <= my_rom(8385); 
 data8 <= my_rom(9740); 
 data9 <= my_rom(11095); 
 data10 <= my_rom(12450);
when "00100000000" => 
 data1 <= my_rom(256); 
 data2 <= my_rom(1611); 
 data3 <= my_rom(2966); 
 data4 <= my_rom(4321); 
 data5 <= my_rom(5676); 
 data6 <= my_rom(7031); 
 data7 <= my_rom(8386); 
 data8 <= my_rom(9741); 
 data9 <= my_rom(11096); 
 data10 <= my_rom(12451);
when "00100000001" => 
 data1 <= my_rom(257); 
 data2 <= my_rom(1612); 
 data3 <= my_rom(2967); 
 data4 <= my_rom(4322); 
 data5 <= my_rom(5677); 
 data6 <= my_rom(7032); 
 data7 <= my_rom(8387); 
 data8 <= my_rom(9742); 
 data9 <= my_rom(11097); 
 data10 <= my_rom(12452);
when "00100000010" => 
 data1 <= my_rom(258); 
 data2 <= my_rom(1613); 
 data3 <= my_rom(2968); 
 data4 <= my_rom(4323); 
 data5 <= my_rom(5678); 
 data6 <= my_rom(7033); 
 data7 <= my_rom(8388); 
 data8 <= my_rom(9743); 
 data9 <= my_rom(11098); 
 data10 <= my_rom(12453);
when "00100000011" => 
 data1 <= my_rom(259); 
 data2 <= my_rom(1614); 
 data3 <= my_rom(2969); 
 data4 <= my_rom(4324); 
 data5 <= my_rom(5679); 
 data6 <= my_rom(7034); 
 data7 <= my_rom(8389); 
 data8 <= my_rom(9744); 
 data9 <= my_rom(11099); 
 data10 <= my_rom(12454);
when "00100000100" => 
 data1 <= my_rom(260); 
 data2 <= my_rom(1615); 
 data3 <= my_rom(2970); 
 data4 <= my_rom(4325); 
 data5 <= my_rom(5680); 
 data6 <= my_rom(7035); 
 data7 <= my_rom(8390); 
 data8 <= my_rom(9745); 
 data9 <= my_rom(11100); 
 data10 <= my_rom(12455);
when "00100000101" => 
 data1 <= my_rom(261); 
 data2 <= my_rom(1616); 
 data3 <= my_rom(2971); 
 data4 <= my_rom(4326); 
 data5 <= my_rom(5681); 
 data6 <= my_rom(7036); 
 data7 <= my_rom(8391); 
 data8 <= my_rom(9746); 
 data9 <= my_rom(11101); 
 data10 <= my_rom(12456);
when "00100000110" => 
 data1 <= my_rom(262); 
 data2 <= my_rom(1617); 
 data3 <= my_rom(2972); 
 data4 <= my_rom(4327); 
 data5 <= my_rom(5682); 
 data6 <= my_rom(7037); 
 data7 <= my_rom(8392); 
 data8 <= my_rom(9747); 
 data9 <= my_rom(11102); 
 data10 <= my_rom(12457);
when "00100000111" => 
 data1 <= my_rom(263); 
 data2 <= my_rom(1618); 
 data3 <= my_rom(2973); 
 data4 <= my_rom(4328); 
 data5 <= my_rom(5683); 
 data6 <= my_rom(7038); 
 data7 <= my_rom(8393); 
 data8 <= my_rom(9748); 
 data9 <= my_rom(11103); 
 data10 <= my_rom(12458);
when "00100001000" => 
 data1 <= my_rom(264); 
 data2 <= my_rom(1619); 
 data3 <= my_rom(2974); 
 data4 <= my_rom(4329); 
 data5 <= my_rom(5684); 
 data6 <= my_rom(7039); 
 data7 <= my_rom(8394); 
 data8 <= my_rom(9749); 
 data9 <= my_rom(11104); 
 data10 <= my_rom(12459);
when "00100001001" => 
 data1 <= my_rom(265); 
 data2 <= my_rom(1620); 
 data3 <= my_rom(2975); 
 data4 <= my_rom(4330); 
 data5 <= my_rom(5685); 
 data6 <= my_rom(7040); 
 data7 <= my_rom(8395); 
 data8 <= my_rom(9750); 
 data9 <= my_rom(11105); 
 data10 <= my_rom(12460);
when "00100001010" => 
 data1 <= my_rom(266); 
 data2 <= my_rom(1621); 
 data3 <= my_rom(2976); 
 data4 <= my_rom(4331); 
 data5 <= my_rom(5686); 
 data6 <= my_rom(7041); 
 data7 <= my_rom(8396); 
 data8 <= my_rom(9751); 
 data9 <= my_rom(11106); 
 data10 <= my_rom(12461);
when "00100001011" => 
 data1 <= my_rom(267); 
 data2 <= my_rom(1622); 
 data3 <= my_rom(2977); 
 data4 <= my_rom(4332); 
 data5 <= my_rom(5687); 
 data6 <= my_rom(7042); 
 data7 <= my_rom(8397); 
 data8 <= my_rom(9752); 
 data9 <= my_rom(11107); 
 data10 <= my_rom(12462);
when "00100001100" => 
 data1 <= my_rom(268); 
 data2 <= my_rom(1623); 
 data3 <= my_rom(2978); 
 data4 <= my_rom(4333); 
 data5 <= my_rom(5688); 
 data6 <= my_rom(7043); 
 data7 <= my_rom(8398); 
 data8 <= my_rom(9753); 
 data9 <= my_rom(11108); 
 data10 <= my_rom(12463);
when "00100001101" => 
 data1 <= my_rom(269); 
 data2 <= my_rom(1624); 
 data3 <= my_rom(2979); 
 data4 <= my_rom(4334); 
 data5 <= my_rom(5689); 
 data6 <= my_rom(7044); 
 data7 <= my_rom(8399); 
 data8 <= my_rom(9754); 
 data9 <= my_rom(11109); 
 data10 <= my_rom(12464);
when "00100001110" => 
 data1 <= my_rom(270); 
 data2 <= my_rom(1625); 
 data3 <= my_rom(2980); 
 data4 <= my_rom(4335); 
 data5 <= my_rom(5690); 
 data6 <= my_rom(7045); 
 data7 <= my_rom(8400); 
 data8 <= my_rom(9755); 
 data9 <= my_rom(11110); 
 data10 <= my_rom(12465);
when "00100001111" => 
 data1 <= my_rom(271); 
 data2 <= my_rom(1626); 
 data3 <= my_rom(2981); 
 data4 <= my_rom(4336); 
 data5 <= my_rom(5691); 
 data6 <= my_rom(7046); 
 data7 <= my_rom(8401); 
 data8 <= my_rom(9756); 
 data9 <= my_rom(11111); 
 data10 <= my_rom(12466);
when "00100010000" => 
 data1 <= my_rom(272); 
 data2 <= my_rom(1627); 
 data3 <= my_rom(2982); 
 data4 <= my_rom(4337); 
 data5 <= my_rom(5692); 
 data6 <= my_rom(7047); 
 data7 <= my_rom(8402); 
 data8 <= my_rom(9757); 
 data9 <= my_rom(11112); 
 data10 <= my_rom(12467);
when "00100010001" => 
 data1 <= my_rom(273); 
 data2 <= my_rom(1628); 
 data3 <= my_rom(2983); 
 data4 <= my_rom(4338); 
 data5 <= my_rom(5693); 
 data6 <= my_rom(7048); 
 data7 <= my_rom(8403); 
 data8 <= my_rom(9758); 
 data9 <= my_rom(11113); 
 data10 <= my_rom(12468);
when "00100010010" => 
 data1 <= my_rom(274); 
 data2 <= my_rom(1629); 
 data3 <= my_rom(2984); 
 data4 <= my_rom(4339); 
 data5 <= my_rom(5694); 
 data6 <= my_rom(7049); 
 data7 <= my_rom(8404); 
 data8 <= my_rom(9759); 
 data9 <= my_rom(11114); 
 data10 <= my_rom(12469);
when "00100010011" => 
 data1 <= my_rom(275); 
 data2 <= my_rom(1630); 
 data3 <= my_rom(2985); 
 data4 <= my_rom(4340); 
 data5 <= my_rom(5695); 
 data6 <= my_rom(7050); 
 data7 <= my_rom(8405); 
 data8 <= my_rom(9760); 
 data9 <= my_rom(11115); 
 data10 <= my_rom(12470);
when "00100010100" => 
 data1 <= my_rom(276); 
 data2 <= my_rom(1631); 
 data3 <= my_rom(2986); 
 data4 <= my_rom(4341); 
 data5 <= my_rom(5696); 
 data6 <= my_rom(7051); 
 data7 <= my_rom(8406); 
 data8 <= my_rom(9761); 
 data9 <= my_rom(11116); 
 data10 <= my_rom(12471);
when "00100010101" => 
 data1 <= my_rom(277); 
 data2 <= my_rom(1632); 
 data3 <= my_rom(2987); 
 data4 <= my_rom(4342); 
 data5 <= my_rom(5697); 
 data6 <= my_rom(7052); 
 data7 <= my_rom(8407); 
 data8 <= my_rom(9762); 
 data9 <= my_rom(11117); 
 data10 <= my_rom(12472);
when "00100010110" => 
 data1 <= my_rom(278); 
 data2 <= my_rom(1633); 
 data3 <= my_rom(2988); 
 data4 <= my_rom(4343); 
 data5 <= my_rom(5698); 
 data6 <= my_rom(7053); 
 data7 <= my_rom(8408); 
 data8 <= my_rom(9763); 
 data9 <= my_rom(11118); 
 data10 <= my_rom(12473);
when "00100010111" => 
 data1 <= my_rom(279); 
 data2 <= my_rom(1634); 
 data3 <= my_rom(2989); 
 data4 <= my_rom(4344); 
 data5 <= my_rom(5699); 
 data6 <= my_rom(7054); 
 data7 <= my_rom(8409); 
 data8 <= my_rom(9764); 
 data9 <= my_rom(11119); 
 data10 <= my_rom(12474);
when "00100011000" => 
 data1 <= my_rom(280); 
 data2 <= my_rom(1635); 
 data3 <= my_rom(2990); 
 data4 <= my_rom(4345); 
 data5 <= my_rom(5700); 
 data6 <= my_rom(7055); 
 data7 <= my_rom(8410); 
 data8 <= my_rom(9765); 
 data9 <= my_rom(11120); 
 data10 <= my_rom(12475);
when "00100011001" => 
 data1 <= my_rom(281); 
 data2 <= my_rom(1636); 
 data3 <= my_rom(2991); 
 data4 <= my_rom(4346); 
 data5 <= my_rom(5701); 
 data6 <= my_rom(7056); 
 data7 <= my_rom(8411); 
 data8 <= my_rom(9766); 
 data9 <= my_rom(11121); 
 data10 <= my_rom(12476);
when "00100011010" => 
 data1 <= my_rom(282); 
 data2 <= my_rom(1637); 
 data3 <= my_rom(2992); 
 data4 <= my_rom(4347); 
 data5 <= my_rom(5702); 
 data6 <= my_rom(7057); 
 data7 <= my_rom(8412); 
 data8 <= my_rom(9767); 
 data9 <= my_rom(11122); 
 data10 <= my_rom(12477);
when "00100011011" => 
 data1 <= my_rom(283); 
 data2 <= my_rom(1638); 
 data3 <= my_rom(2993); 
 data4 <= my_rom(4348); 
 data5 <= my_rom(5703); 
 data6 <= my_rom(7058); 
 data7 <= my_rom(8413); 
 data8 <= my_rom(9768); 
 data9 <= my_rom(11123); 
 data10 <= my_rom(12478);
when "00100011100" => 
 data1 <= my_rom(284); 
 data2 <= my_rom(1639); 
 data3 <= my_rom(2994); 
 data4 <= my_rom(4349); 
 data5 <= my_rom(5704); 
 data6 <= my_rom(7059); 
 data7 <= my_rom(8414); 
 data8 <= my_rom(9769); 
 data9 <= my_rom(11124); 
 data10 <= my_rom(12479);
when "00100011101" => 
 data1 <= my_rom(285); 
 data2 <= my_rom(1640); 
 data3 <= my_rom(2995); 
 data4 <= my_rom(4350); 
 data5 <= my_rom(5705); 
 data6 <= my_rom(7060); 
 data7 <= my_rom(8415); 
 data8 <= my_rom(9770); 
 data9 <= my_rom(11125); 
 data10 <= my_rom(12480);
when "00100011110" => 
 data1 <= my_rom(286); 
 data2 <= my_rom(1641); 
 data3 <= my_rom(2996); 
 data4 <= my_rom(4351); 
 data5 <= my_rom(5706); 
 data6 <= my_rom(7061); 
 data7 <= my_rom(8416); 
 data8 <= my_rom(9771); 
 data9 <= my_rom(11126); 
 data10 <= my_rom(12481);
when "00100011111" => 
 data1 <= my_rom(287); 
 data2 <= my_rom(1642); 
 data3 <= my_rom(2997); 
 data4 <= my_rom(4352); 
 data5 <= my_rom(5707); 
 data6 <= my_rom(7062); 
 data7 <= my_rom(8417); 
 data8 <= my_rom(9772); 
 data9 <= my_rom(11127); 
 data10 <= my_rom(12482);
when "00100100000" => 
 data1 <= my_rom(288); 
 data2 <= my_rom(1643); 
 data3 <= my_rom(2998); 
 data4 <= my_rom(4353); 
 data5 <= my_rom(5708); 
 data6 <= my_rom(7063); 
 data7 <= my_rom(8418); 
 data8 <= my_rom(9773); 
 data9 <= my_rom(11128); 
 data10 <= my_rom(12483);
when "00100100001" => 
 data1 <= my_rom(289); 
 data2 <= my_rom(1644); 
 data3 <= my_rom(2999); 
 data4 <= my_rom(4354); 
 data5 <= my_rom(5709); 
 data6 <= my_rom(7064); 
 data7 <= my_rom(8419); 
 data8 <= my_rom(9774); 
 data9 <= my_rom(11129); 
 data10 <= my_rom(12484);
when "00100100010" => 
 data1 <= my_rom(290); 
 data2 <= my_rom(1645); 
 data3 <= my_rom(3000); 
 data4 <= my_rom(4355); 
 data5 <= my_rom(5710); 
 data6 <= my_rom(7065); 
 data7 <= my_rom(8420); 
 data8 <= my_rom(9775); 
 data9 <= my_rom(11130); 
 data10 <= my_rom(12485);
when "00100100011" => 
 data1 <= my_rom(291); 
 data2 <= my_rom(1646); 
 data3 <= my_rom(3001); 
 data4 <= my_rom(4356); 
 data5 <= my_rom(5711); 
 data6 <= my_rom(7066); 
 data7 <= my_rom(8421); 
 data8 <= my_rom(9776); 
 data9 <= my_rom(11131); 
 data10 <= my_rom(12486);
when "00100100100" => 
 data1 <= my_rom(292); 
 data2 <= my_rom(1647); 
 data3 <= my_rom(3002); 
 data4 <= my_rom(4357); 
 data5 <= my_rom(5712); 
 data6 <= my_rom(7067); 
 data7 <= my_rom(8422); 
 data8 <= my_rom(9777); 
 data9 <= my_rom(11132); 
 data10 <= my_rom(12487);
when "00100100101" => 
 data1 <= my_rom(293); 
 data2 <= my_rom(1648); 
 data3 <= my_rom(3003); 
 data4 <= my_rom(4358); 
 data5 <= my_rom(5713); 
 data6 <= my_rom(7068); 
 data7 <= my_rom(8423); 
 data8 <= my_rom(9778); 
 data9 <= my_rom(11133); 
 data10 <= my_rom(12488);
when "00100100110" => 
 data1 <= my_rom(294); 
 data2 <= my_rom(1649); 
 data3 <= my_rom(3004); 
 data4 <= my_rom(4359); 
 data5 <= my_rom(5714); 
 data6 <= my_rom(7069); 
 data7 <= my_rom(8424); 
 data8 <= my_rom(9779); 
 data9 <= my_rom(11134); 
 data10 <= my_rom(12489);
when "00100100111" => 
 data1 <= my_rom(295); 
 data2 <= my_rom(1650); 
 data3 <= my_rom(3005); 
 data4 <= my_rom(4360); 
 data5 <= my_rom(5715); 
 data6 <= my_rom(7070); 
 data7 <= my_rom(8425); 
 data8 <= my_rom(9780); 
 data9 <= my_rom(11135); 
 data10 <= my_rom(12490);
when "00100101000" => 
 data1 <= my_rom(296); 
 data2 <= my_rom(1651); 
 data3 <= my_rom(3006); 
 data4 <= my_rom(4361); 
 data5 <= my_rom(5716); 
 data6 <= my_rom(7071); 
 data7 <= my_rom(8426); 
 data8 <= my_rom(9781); 
 data9 <= my_rom(11136); 
 data10 <= my_rom(12491);
when "00100101001" => 
 data1 <= my_rom(297); 
 data2 <= my_rom(1652); 
 data3 <= my_rom(3007); 
 data4 <= my_rom(4362); 
 data5 <= my_rom(5717); 
 data6 <= my_rom(7072); 
 data7 <= my_rom(8427); 
 data8 <= my_rom(9782); 
 data9 <= my_rom(11137); 
 data10 <= my_rom(12492);
when "00100101010" => 
 data1 <= my_rom(298); 
 data2 <= my_rom(1653); 
 data3 <= my_rom(3008); 
 data4 <= my_rom(4363); 
 data5 <= my_rom(5718); 
 data6 <= my_rom(7073); 
 data7 <= my_rom(8428); 
 data8 <= my_rom(9783); 
 data9 <= my_rom(11138); 
 data10 <= my_rom(12493);
when "00100101011" => 
 data1 <= my_rom(299); 
 data2 <= my_rom(1654); 
 data3 <= my_rom(3009); 
 data4 <= my_rom(4364); 
 data5 <= my_rom(5719); 
 data6 <= my_rom(7074); 
 data7 <= my_rom(8429); 
 data8 <= my_rom(9784); 
 data9 <= my_rom(11139); 
 data10 <= my_rom(12494);
when "00100101100" => 
 data1 <= my_rom(300); 
 data2 <= my_rom(1655); 
 data3 <= my_rom(3010); 
 data4 <= my_rom(4365); 
 data5 <= my_rom(5720); 
 data6 <= my_rom(7075); 
 data7 <= my_rom(8430); 
 data8 <= my_rom(9785); 
 data9 <= my_rom(11140); 
 data10 <= my_rom(12495);
when "00100101101" => 
 data1 <= my_rom(301); 
 data2 <= my_rom(1656); 
 data3 <= my_rom(3011); 
 data4 <= my_rom(4366); 
 data5 <= my_rom(5721); 
 data6 <= my_rom(7076); 
 data7 <= my_rom(8431); 
 data8 <= my_rom(9786); 
 data9 <= my_rom(11141); 
 data10 <= my_rom(12496);
when "00100101110" => 
 data1 <= my_rom(302); 
 data2 <= my_rom(1657); 
 data3 <= my_rom(3012); 
 data4 <= my_rom(4367); 
 data5 <= my_rom(5722); 
 data6 <= my_rom(7077); 
 data7 <= my_rom(8432); 
 data8 <= my_rom(9787); 
 data9 <= my_rom(11142); 
 data10 <= my_rom(12497);
when "00100101111" => 
 data1 <= my_rom(303); 
 data2 <= my_rom(1658); 
 data3 <= my_rom(3013); 
 data4 <= my_rom(4368); 
 data5 <= my_rom(5723); 
 data6 <= my_rom(7078); 
 data7 <= my_rom(8433); 
 data8 <= my_rom(9788); 
 data9 <= my_rom(11143); 
 data10 <= my_rom(12498);
when "00100110000" => 
 data1 <= my_rom(304); 
 data2 <= my_rom(1659); 
 data3 <= my_rom(3014); 
 data4 <= my_rom(4369); 
 data5 <= my_rom(5724); 
 data6 <= my_rom(7079); 
 data7 <= my_rom(8434); 
 data8 <= my_rom(9789); 
 data9 <= my_rom(11144); 
 data10 <= my_rom(12499);
when "00100110001" => 
 data1 <= my_rom(305); 
 data2 <= my_rom(1660); 
 data3 <= my_rom(3015); 
 data4 <= my_rom(4370); 
 data5 <= my_rom(5725); 
 data6 <= my_rom(7080); 
 data7 <= my_rom(8435); 
 data8 <= my_rom(9790); 
 data9 <= my_rom(11145); 
 data10 <= my_rom(12500);
when "00100110010" => 
 data1 <= my_rom(306); 
 data2 <= my_rom(1661); 
 data3 <= my_rom(3016); 
 data4 <= my_rom(4371); 
 data5 <= my_rom(5726); 
 data6 <= my_rom(7081); 
 data7 <= my_rom(8436); 
 data8 <= my_rom(9791); 
 data9 <= my_rom(11146); 
 data10 <= my_rom(12501);
when "00100110011" => 
 data1 <= my_rom(307); 
 data2 <= my_rom(1662); 
 data3 <= my_rom(3017); 
 data4 <= my_rom(4372); 
 data5 <= my_rom(5727); 
 data6 <= my_rom(7082); 
 data7 <= my_rom(8437); 
 data8 <= my_rom(9792); 
 data9 <= my_rom(11147); 
 data10 <= my_rom(12502);
when "00100110100" => 
 data1 <= my_rom(308); 
 data2 <= my_rom(1663); 
 data3 <= my_rom(3018); 
 data4 <= my_rom(4373); 
 data5 <= my_rom(5728); 
 data6 <= my_rom(7083); 
 data7 <= my_rom(8438); 
 data8 <= my_rom(9793); 
 data9 <= my_rom(11148); 
 data10 <= my_rom(12503);
when "00100110101" => 
 data1 <= my_rom(309); 
 data2 <= my_rom(1664); 
 data3 <= my_rom(3019); 
 data4 <= my_rom(4374); 
 data5 <= my_rom(5729); 
 data6 <= my_rom(7084); 
 data7 <= my_rom(8439); 
 data8 <= my_rom(9794); 
 data9 <= my_rom(11149); 
 data10 <= my_rom(12504);
when "00100110110" => 
 data1 <= my_rom(310); 
 data2 <= my_rom(1665); 
 data3 <= my_rom(3020); 
 data4 <= my_rom(4375); 
 data5 <= my_rom(5730); 
 data6 <= my_rom(7085); 
 data7 <= my_rom(8440); 
 data8 <= my_rom(9795); 
 data9 <= my_rom(11150); 
 data10 <= my_rom(12505);
when "00100110111" => 
 data1 <= my_rom(311); 
 data2 <= my_rom(1666); 
 data3 <= my_rom(3021); 
 data4 <= my_rom(4376); 
 data5 <= my_rom(5731); 
 data6 <= my_rom(7086); 
 data7 <= my_rom(8441); 
 data8 <= my_rom(9796); 
 data9 <= my_rom(11151); 
 data10 <= my_rom(12506);
when "00100111000" => 
 data1 <= my_rom(312); 
 data2 <= my_rom(1667); 
 data3 <= my_rom(3022); 
 data4 <= my_rom(4377); 
 data5 <= my_rom(5732); 
 data6 <= my_rom(7087); 
 data7 <= my_rom(8442); 
 data8 <= my_rom(9797); 
 data9 <= my_rom(11152); 
 data10 <= my_rom(12507);
when "00100111001" => 
 data1 <= my_rom(313); 
 data2 <= my_rom(1668); 
 data3 <= my_rom(3023); 
 data4 <= my_rom(4378); 
 data5 <= my_rom(5733); 
 data6 <= my_rom(7088); 
 data7 <= my_rom(8443); 
 data8 <= my_rom(9798); 
 data9 <= my_rom(11153); 
 data10 <= my_rom(12508);
when "00100111010" => 
 data1 <= my_rom(314); 
 data2 <= my_rom(1669); 
 data3 <= my_rom(3024); 
 data4 <= my_rom(4379); 
 data5 <= my_rom(5734); 
 data6 <= my_rom(7089); 
 data7 <= my_rom(8444); 
 data8 <= my_rom(9799); 
 data9 <= my_rom(11154); 
 data10 <= my_rom(12509);
when "00100111011" => 
 data1 <= my_rom(315); 
 data2 <= my_rom(1670); 
 data3 <= my_rom(3025); 
 data4 <= my_rom(4380); 
 data5 <= my_rom(5735); 
 data6 <= my_rom(7090); 
 data7 <= my_rom(8445); 
 data8 <= my_rom(9800); 
 data9 <= my_rom(11155); 
 data10 <= my_rom(12510);
when "00100111100" => 
 data1 <= my_rom(316); 
 data2 <= my_rom(1671); 
 data3 <= my_rom(3026); 
 data4 <= my_rom(4381); 
 data5 <= my_rom(5736); 
 data6 <= my_rom(7091); 
 data7 <= my_rom(8446); 
 data8 <= my_rom(9801); 
 data9 <= my_rom(11156); 
 data10 <= my_rom(12511);
when "00100111101" => 
 data1 <= my_rom(317); 
 data2 <= my_rom(1672); 
 data3 <= my_rom(3027); 
 data4 <= my_rom(4382); 
 data5 <= my_rom(5737); 
 data6 <= my_rom(7092); 
 data7 <= my_rom(8447); 
 data8 <= my_rom(9802); 
 data9 <= my_rom(11157); 
 data10 <= my_rom(12512);
when "00100111110" => 
 data1 <= my_rom(318); 
 data2 <= my_rom(1673); 
 data3 <= my_rom(3028); 
 data4 <= my_rom(4383); 
 data5 <= my_rom(5738); 
 data6 <= my_rom(7093); 
 data7 <= my_rom(8448); 
 data8 <= my_rom(9803); 
 data9 <= my_rom(11158); 
 data10 <= my_rom(12513);
when "00100111111" => 
 data1 <= my_rom(319); 
 data2 <= my_rom(1674); 
 data3 <= my_rom(3029); 
 data4 <= my_rom(4384); 
 data5 <= my_rom(5739); 
 data6 <= my_rom(7094); 
 data7 <= my_rom(8449); 
 data8 <= my_rom(9804); 
 data9 <= my_rom(11159); 
 data10 <= my_rom(12514);
when "00101000000" => 
 data1 <= my_rom(320); 
 data2 <= my_rom(1675); 
 data3 <= my_rom(3030); 
 data4 <= my_rom(4385); 
 data5 <= my_rom(5740); 
 data6 <= my_rom(7095); 
 data7 <= my_rom(8450); 
 data8 <= my_rom(9805); 
 data9 <= my_rom(11160); 
 data10 <= my_rom(12515);
when "00101000001" => 
 data1 <= my_rom(321); 
 data2 <= my_rom(1676); 
 data3 <= my_rom(3031); 
 data4 <= my_rom(4386); 
 data5 <= my_rom(5741); 
 data6 <= my_rom(7096); 
 data7 <= my_rom(8451); 
 data8 <= my_rom(9806); 
 data9 <= my_rom(11161); 
 data10 <= my_rom(12516);
when "00101000010" => 
 data1 <= my_rom(322); 
 data2 <= my_rom(1677); 
 data3 <= my_rom(3032); 
 data4 <= my_rom(4387); 
 data5 <= my_rom(5742); 
 data6 <= my_rom(7097); 
 data7 <= my_rom(8452); 
 data8 <= my_rom(9807); 
 data9 <= my_rom(11162); 
 data10 <= my_rom(12517);
when "00101000011" => 
 data1 <= my_rom(323); 
 data2 <= my_rom(1678); 
 data3 <= my_rom(3033); 
 data4 <= my_rom(4388); 
 data5 <= my_rom(5743); 
 data6 <= my_rom(7098); 
 data7 <= my_rom(8453); 
 data8 <= my_rom(9808); 
 data9 <= my_rom(11163); 
 data10 <= my_rom(12518);
when "00101000100" => 
 data1 <= my_rom(324); 
 data2 <= my_rom(1679); 
 data3 <= my_rom(3034); 
 data4 <= my_rom(4389); 
 data5 <= my_rom(5744); 
 data6 <= my_rom(7099); 
 data7 <= my_rom(8454); 
 data8 <= my_rom(9809); 
 data9 <= my_rom(11164); 
 data10 <= my_rom(12519);
when "00101000101" => 
 data1 <= my_rom(325); 
 data2 <= my_rom(1680); 
 data3 <= my_rom(3035); 
 data4 <= my_rom(4390); 
 data5 <= my_rom(5745); 
 data6 <= my_rom(7100); 
 data7 <= my_rom(8455); 
 data8 <= my_rom(9810); 
 data9 <= my_rom(11165); 
 data10 <= my_rom(12520);
when "00101000110" => 
 data1 <= my_rom(326); 
 data2 <= my_rom(1681); 
 data3 <= my_rom(3036); 
 data4 <= my_rom(4391); 
 data5 <= my_rom(5746); 
 data6 <= my_rom(7101); 
 data7 <= my_rom(8456); 
 data8 <= my_rom(9811); 
 data9 <= my_rom(11166); 
 data10 <= my_rom(12521);
when "00101000111" => 
 data1 <= my_rom(327); 
 data2 <= my_rom(1682); 
 data3 <= my_rom(3037); 
 data4 <= my_rom(4392); 
 data5 <= my_rom(5747); 
 data6 <= my_rom(7102); 
 data7 <= my_rom(8457); 
 data8 <= my_rom(9812); 
 data9 <= my_rom(11167); 
 data10 <= my_rom(12522);
when "00101001000" => 
 data1 <= my_rom(328); 
 data2 <= my_rom(1683); 
 data3 <= my_rom(3038); 
 data4 <= my_rom(4393); 
 data5 <= my_rom(5748); 
 data6 <= my_rom(7103); 
 data7 <= my_rom(8458); 
 data8 <= my_rom(9813); 
 data9 <= my_rom(11168); 
 data10 <= my_rom(12523);
when "00101001001" => 
 data1 <= my_rom(329); 
 data2 <= my_rom(1684); 
 data3 <= my_rom(3039); 
 data4 <= my_rom(4394); 
 data5 <= my_rom(5749); 
 data6 <= my_rom(7104); 
 data7 <= my_rom(8459); 
 data8 <= my_rom(9814); 
 data9 <= my_rom(11169); 
 data10 <= my_rom(12524);
when "00101001010" => 
 data1 <= my_rom(330); 
 data2 <= my_rom(1685); 
 data3 <= my_rom(3040); 
 data4 <= my_rom(4395); 
 data5 <= my_rom(5750); 
 data6 <= my_rom(7105); 
 data7 <= my_rom(8460); 
 data8 <= my_rom(9815); 
 data9 <= my_rom(11170); 
 data10 <= my_rom(12525);
when "00101001011" => 
 data1 <= my_rom(331); 
 data2 <= my_rom(1686); 
 data3 <= my_rom(3041); 
 data4 <= my_rom(4396); 
 data5 <= my_rom(5751); 
 data6 <= my_rom(7106); 
 data7 <= my_rom(8461); 
 data8 <= my_rom(9816); 
 data9 <= my_rom(11171); 
 data10 <= my_rom(12526);
when "00101001100" => 
 data1 <= my_rom(332); 
 data2 <= my_rom(1687); 
 data3 <= my_rom(3042); 
 data4 <= my_rom(4397); 
 data5 <= my_rom(5752); 
 data6 <= my_rom(7107); 
 data7 <= my_rom(8462); 
 data8 <= my_rom(9817); 
 data9 <= my_rom(11172); 
 data10 <= my_rom(12527);
when "00101001101" => 
 data1 <= my_rom(333); 
 data2 <= my_rom(1688); 
 data3 <= my_rom(3043); 
 data4 <= my_rom(4398); 
 data5 <= my_rom(5753); 
 data6 <= my_rom(7108); 
 data7 <= my_rom(8463); 
 data8 <= my_rom(9818); 
 data9 <= my_rom(11173); 
 data10 <= my_rom(12528);
when "00101001110" => 
 data1 <= my_rom(334); 
 data2 <= my_rom(1689); 
 data3 <= my_rom(3044); 
 data4 <= my_rom(4399); 
 data5 <= my_rom(5754); 
 data6 <= my_rom(7109); 
 data7 <= my_rom(8464); 
 data8 <= my_rom(9819); 
 data9 <= my_rom(11174); 
 data10 <= my_rom(12529);
when "00101001111" => 
 data1 <= my_rom(335); 
 data2 <= my_rom(1690); 
 data3 <= my_rom(3045); 
 data4 <= my_rom(4400); 
 data5 <= my_rom(5755); 
 data6 <= my_rom(7110); 
 data7 <= my_rom(8465); 
 data8 <= my_rom(9820); 
 data9 <= my_rom(11175); 
 data10 <= my_rom(12530);
when "00101010000" => 
 data1 <= my_rom(336); 
 data2 <= my_rom(1691); 
 data3 <= my_rom(3046); 
 data4 <= my_rom(4401); 
 data5 <= my_rom(5756); 
 data6 <= my_rom(7111); 
 data7 <= my_rom(8466); 
 data8 <= my_rom(9821); 
 data9 <= my_rom(11176); 
 data10 <= my_rom(12531);
when "00101010001" => 
 data1 <= my_rom(337); 
 data2 <= my_rom(1692); 
 data3 <= my_rom(3047); 
 data4 <= my_rom(4402); 
 data5 <= my_rom(5757); 
 data6 <= my_rom(7112); 
 data7 <= my_rom(8467); 
 data8 <= my_rom(9822); 
 data9 <= my_rom(11177); 
 data10 <= my_rom(12532);
when "00101010010" => 
 data1 <= my_rom(338); 
 data2 <= my_rom(1693); 
 data3 <= my_rom(3048); 
 data4 <= my_rom(4403); 
 data5 <= my_rom(5758); 
 data6 <= my_rom(7113); 
 data7 <= my_rom(8468); 
 data8 <= my_rom(9823); 
 data9 <= my_rom(11178); 
 data10 <= my_rom(12533);
when "00101010011" => 
 data1 <= my_rom(339); 
 data2 <= my_rom(1694); 
 data3 <= my_rom(3049); 
 data4 <= my_rom(4404); 
 data5 <= my_rom(5759); 
 data6 <= my_rom(7114); 
 data7 <= my_rom(8469); 
 data8 <= my_rom(9824); 
 data9 <= my_rom(11179); 
 data10 <= my_rom(12534);
when "00101010100" => 
 data1 <= my_rom(340); 
 data2 <= my_rom(1695); 
 data3 <= my_rom(3050); 
 data4 <= my_rom(4405); 
 data5 <= my_rom(5760); 
 data6 <= my_rom(7115); 
 data7 <= my_rom(8470); 
 data8 <= my_rom(9825); 
 data9 <= my_rom(11180); 
 data10 <= my_rom(12535);
when "00101010101" => 
 data1 <= my_rom(341); 
 data2 <= my_rom(1696); 
 data3 <= my_rom(3051); 
 data4 <= my_rom(4406); 
 data5 <= my_rom(5761); 
 data6 <= my_rom(7116); 
 data7 <= my_rom(8471); 
 data8 <= my_rom(9826); 
 data9 <= my_rom(11181); 
 data10 <= my_rom(12536);
when "00101010110" => 
 data1 <= my_rom(342); 
 data2 <= my_rom(1697); 
 data3 <= my_rom(3052); 
 data4 <= my_rom(4407); 
 data5 <= my_rom(5762); 
 data6 <= my_rom(7117); 
 data7 <= my_rom(8472); 
 data8 <= my_rom(9827); 
 data9 <= my_rom(11182); 
 data10 <= my_rom(12537);
when "00101010111" => 
 data1 <= my_rom(343); 
 data2 <= my_rom(1698); 
 data3 <= my_rom(3053); 
 data4 <= my_rom(4408); 
 data5 <= my_rom(5763); 
 data6 <= my_rom(7118); 
 data7 <= my_rom(8473); 
 data8 <= my_rom(9828); 
 data9 <= my_rom(11183); 
 data10 <= my_rom(12538);
when "00101011000" => 
 data1 <= my_rom(344); 
 data2 <= my_rom(1699); 
 data3 <= my_rom(3054); 
 data4 <= my_rom(4409); 
 data5 <= my_rom(5764); 
 data6 <= my_rom(7119); 
 data7 <= my_rom(8474); 
 data8 <= my_rom(9829); 
 data9 <= my_rom(11184); 
 data10 <= my_rom(12539);
when "00101011001" => 
 data1 <= my_rom(345); 
 data2 <= my_rom(1700); 
 data3 <= my_rom(3055); 
 data4 <= my_rom(4410); 
 data5 <= my_rom(5765); 
 data6 <= my_rom(7120); 
 data7 <= my_rom(8475); 
 data8 <= my_rom(9830); 
 data9 <= my_rom(11185); 
 data10 <= my_rom(12540);
when "00101011010" => 
 data1 <= my_rom(346); 
 data2 <= my_rom(1701); 
 data3 <= my_rom(3056); 
 data4 <= my_rom(4411); 
 data5 <= my_rom(5766); 
 data6 <= my_rom(7121); 
 data7 <= my_rom(8476); 
 data8 <= my_rom(9831); 
 data9 <= my_rom(11186); 
 data10 <= my_rom(12541);
when "00101011011" => 
 data1 <= my_rom(347); 
 data2 <= my_rom(1702); 
 data3 <= my_rom(3057); 
 data4 <= my_rom(4412); 
 data5 <= my_rom(5767); 
 data6 <= my_rom(7122); 
 data7 <= my_rom(8477); 
 data8 <= my_rom(9832); 
 data9 <= my_rom(11187); 
 data10 <= my_rom(12542);
when "00101011100" => 
 data1 <= my_rom(348); 
 data2 <= my_rom(1703); 
 data3 <= my_rom(3058); 
 data4 <= my_rom(4413); 
 data5 <= my_rom(5768); 
 data6 <= my_rom(7123); 
 data7 <= my_rom(8478); 
 data8 <= my_rom(9833); 
 data9 <= my_rom(11188); 
 data10 <= my_rom(12543);
when "00101011101" => 
 data1 <= my_rom(349); 
 data2 <= my_rom(1704); 
 data3 <= my_rom(3059); 
 data4 <= my_rom(4414); 
 data5 <= my_rom(5769); 
 data6 <= my_rom(7124); 
 data7 <= my_rom(8479); 
 data8 <= my_rom(9834); 
 data9 <= my_rom(11189); 
 data10 <= my_rom(12544);
when "00101011110" => 
 data1 <= my_rom(350); 
 data2 <= my_rom(1705); 
 data3 <= my_rom(3060); 
 data4 <= my_rom(4415); 
 data5 <= my_rom(5770); 
 data6 <= my_rom(7125); 
 data7 <= my_rom(8480); 
 data8 <= my_rom(9835); 
 data9 <= my_rom(11190); 
 data10 <= my_rom(12545);
when "00101011111" => 
 data1 <= my_rom(351); 
 data2 <= my_rom(1706); 
 data3 <= my_rom(3061); 
 data4 <= my_rom(4416); 
 data5 <= my_rom(5771); 
 data6 <= my_rom(7126); 
 data7 <= my_rom(8481); 
 data8 <= my_rom(9836); 
 data9 <= my_rom(11191); 
 data10 <= my_rom(12546);
when "00101100000" => 
 data1 <= my_rom(352); 
 data2 <= my_rom(1707); 
 data3 <= my_rom(3062); 
 data4 <= my_rom(4417); 
 data5 <= my_rom(5772); 
 data6 <= my_rom(7127); 
 data7 <= my_rom(8482); 
 data8 <= my_rom(9837); 
 data9 <= my_rom(11192); 
 data10 <= my_rom(12547);
when "00101100001" => 
 data1 <= my_rom(353); 
 data2 <= my_rom(1708); 
 data3 <= my_rom(3063); 
 data4 <= my_rom(4418); 
 data5 <= my_rom(5773); 
 data6 <= my_rom(7128); 
 data7 <= my_rom(8483); 
 data8 <= my_rom(9838); 
 data9 <= my_rom(11193); 
 data10 <= my_rom(12548);
when "00101100010" => 
 data1 <= my_rom(354); 
 data2 <= my_rom(1709); 
 data3 <= my_rom(3064); 
 data4 <= my_rom(4419); 
 data5 <= my_rom(5774); 
 data6 <= my_rom(7129); 
 data7 <= my_rom(8484); 
 data8 <= my_rom(9839); 
 data9 <= my_rom(11194); 
 data10 <= my_rom(12549);
when "00101100011" => 
 data1 <= my_rom(355); 
 data2 <= my_rom(1710); 
 data3 <= my_rom(3065); 
 data4 <= my_rom(4420); 
 data5 <= my_rom(5775); 
 data6 <= my_rom(7130); 
 data7 <= my_rom(8485); 
 data8 <= my_rom(9840); 
 data9 <= my_rom(11195); 
 data10 <= my_rom(12550);
when "00101100100" => 
 data1 <= my_rom(356); 
 data2 <= my_rom(1711); 
 data3 <= my_rom(3066); 
 data4 <= my_rom(4421); 
 data5 <= my_rom(5776); 
 data6 <= my_rom(7131); 
 data7 <= my_rom(8486); 
 data8 <= my_rom(9841); 
 data9 <= my_rom(11196); 
 data10 <= my_rom(12551);
when "00101100101" => 
 data1 <= my_rom(357); 
 data2 <= my_rom(1712); 
 data3 <= my_rom(3067); 
 data4 <= my_rom(4422); 
 data5 <= my_rom(5777); 
 data6 <= my_rom(7132); 
 data7 <= my_rom(8487); 
 data8 <= my_rom(9842); 
 data9 <= my_rom(11197); 
 data10 <= my_rom(12552);
when "00101100110" => 
 data1 <= my_rom(358); 
 data2 <= my_rom(1713); 
 data3 <= my_rom(3068); 
 data4 <= my_rom(4423); 
 data5 <= my_rom(5778); 
 data6 <= my_rom(7133); 
 data7 <= my_rom(8488); 
 data8 <= my_rom(9843); 
 data9 <= my_rom(11198); 
 data10 <= my_rom(12553);
when "00101100111" => 
 data1 <= my_rom(359); 
 data2 <= my_rom(1714); 
 data3 <= my_rom(3069); 
 data4 <= my_rom(4424); 
 data5 <= my_rom(5779); 
 data6 <= my_rom(7134); 
 data7 <= my_rom(8489); 
 data8 <= my_rom(9844); 
 data9 <= my_rom(11199); 
 data10 <= my_rom(12554);
when "00101101000" => 
 data1 <= my_rom(360); 
 data2 <= my_rom(1715); 
 data3 <= my_rom(3070); 
 data4 <= my_rom(4425); 
 data5 <= my_rom(5780); 
 data6 <= my_rom(7135); 
 data7 <= my_rom(8490); 
 data8 <= my_rom(9845); 
 data9 <= my_rom(11200); 
 data10 <= my_rom(12555);
when "00101101001" => 
 data1 <= my_rom(361); 
 data2 <= my_rom(1716); 
 data3 <= my_rom(3071); 
 data4 <= my_rom(4426); 
 data5 <= my_rom(5781); 
 data6 <= my_rom(7136); 
 data7 <= my_rom(8491); 
 data8 <= my_rom(9846); 
 data9 <= my_rom(11201); 
 data10 <= my_rom(12556);
when "00101101010" => 
 data1 <= my_rom(362); 
 data2 <= my_rom(1717); 
 data3 <= my_rom(3072); 
 data4 <= my_rom(4427); 
 data5 <= my_rom(5782); 
 data6 <= my_rom(7137); 
 data7 <= my_rom(8492); 
 data8 <= my_rom(9847); 
 data9 <= my_rom(11202); 
 data10 <= my_rom(12557);
when "00101101011" => 
 data1 <= my_rom(363); 
 data2 <= my_rom(1718); 
 data3 <= my_rom(3073); 
 data4 <= my_rom(4428); 
 data5 <= my_rom(5783); 
 data6 <= my_rom(7138); 
 data7 <= my_rom(8493); 
 data8 <= my_rom(9848); 
 data9 <= my_rom(11203); 
 data10 <= my_rom(12558);
when "00101101100" => 
 data1 <= my_rom(364); 
 data2 <= my_rom(1719); 
 data3 <= my_rom(3074); 
 data4 <= my_rom(4429); 
 data5 <= my_rom(5784); 
 data6 <= my_rom(7139); 
 data7 <= my_rom(8494); 
 data8 <= my_rom(9849); 
 data9 <= my_rom(11204); 
 data10 <= my_rom(12559);
when "00101101101" => 
 data1 <= my_rom(365); 
 data2 <= my_rom(1720); 
 data3 <= my_rom(3075); 
 data4 <= my_rom(4430); 
 data5 <= my_rom(5785); 
 data6 <= my_rom(7140); 
 data7 <= my_rom(8495); 
 data8 <= my_rom(9850); 
 data9 <= my_rom(11205); 
 data10 <= my_rom(12560);
when "00101101110" => 
 data1 <= my_rom(366); 
 data2 <= my_rom(1721); 
 data3 <= my_rom(3076); 
 data4 <= my_rom(4431); 
 data5 <= my_rom(5786); 
 data6 <= my_rom(7141); 
 data7 <= my_rom(8496); 
 data8 <= my_rom(9851); 
 data9 <= my_rom(11206); 
 data10 <= my_rom(12561);
when "00101101111" => 
 data1 <= my_rom(367); 
 data2 <= my_rom(1722); 
 data3 <= my_rom(3077); 
 data4 <= my_rom(4432); 
 data5 <= my_rom(5787); 
 data6 <= my_rom(7142); 
 data7 <= my_rom(8497); 
 data8 <= my_rom(9852); 
 data9 <= my_rom(11207); 
 data10 <= my_rom(12562);
when "00101110000" => 
 data1 <= my_rom(368); 
 data2 <= my_rom(1723); 
 data3 <= my_rom(3078); 
 data4 <= my_rom(4433); 
 data5 <= my_rom(5788); 
 data6 <= my_rom(7143); 
 data7 <= my_rom(8498); 
 data8 <= my_rom(9853); 
 data9 <= my_rom(11208); 
 data10 <= my_rom(12563);
when "00101110001" => 
 data1 <= my_rom(369); 
 data2 <= my_rom(1724); 
 data3 <= my_rom(3079); 
 data4 <= my_rom(4434); 
 data5 <= my_rom(5789); 
 data6 <= my_rom(7144); 
 data7 <= my_rom(8499); 
 data8 <= my_rom(9854); 
 data9 <= my_rom(11209); 
 data10 <= my_rom(12564);
when "00101110010" => 
 data1 <= my_rom(370); 
 data2 <= my_rom(1725); 
 data3 <= my_rom(3080); 
 data4 <= my_rom(4435); 
 data5 <= my_rom(5790); 
 data6 <= my_rom(7145); 
 data7 <= my_rom(8500); 
 data8 <= my_rom(9855); 
 data9 <= my_rom(11210); 
 data10 <= my_rom(12565);
when "00101110011" => 
 data1 <= my_rom(371); 
 data2 <= my_rom(1726); 
 data3 <= my_rom(3081); 
 data4 <= my_rom(4436); 
 data5 <= my_rom(5791); 
 data6 <= my_rom(7146); 
 data7 <= my_rom(8501); 
 data8 <= my_rom(9856); 
 data9 <= my_rom(11211); 
 data10 <= my_rom(12566);
when "00101110100" => 
 data1 <= my_rom(372); 
 data2 <= my_rom(1727); 
 data3 <= my_rom(3082); 
 data4 <= my_rom(4437); 
 data5 <= my_rom(5792); 
 data6 <= my_rom(7147); 
 data7 <= my_rom(8502); 
 data8 <= my_rom(9857); 
 data9 <= my_rom(11212); 
 data10 <= my_rom(12567);
when "00101110101" => 
 data1 <= my_rom(373); 
 data2 <= my_rom(1728); 
 data3 <= my_rom(3083); 
 data4 <= my_rom(4438); 
 data5 <= my_rom(5793); 
 data6 <= my_rom(7148); 
 data7 <= my_rom(8503); 
 data8 <= my_rom(9858); 
 data9 <= my_rom(11213); 
 data10 <= my_rom(12568);
when "00101110110" => 
 data1 <= my_rom(374); 
 data2 <= my_rom(1729); 
 data3 <= my_rom(3084); 
 data4 <= my_rom(4439); 
 data5 <= my_rom(5794); 
 data6 <= my_rom(7149); 
 data7 <= my_rom(8504); 
 data8 <= my_rom(9859); 
 data9 <= my_rom(11214); 
 data10 <= my_rom(12569);
when "00101110111" => 
 data1 <= my_rom(375); 
 data2 <= my_rom(1730); 
 data3 <= my_rom(3085); 
 data4 <= my_rom(4440); 
 data5 <= my_rom(5795); 
 data6 <= my_rom(7150); 
 data7 <= my_rom(8505); 
 data8 <= my_rom(9860); 
 data9 <= my_rom(11215); 
 data10 <= my_rom(12570);
when "00101111000" => 
 data1 <= my_rom(376); 
 data2 <= my_rom(1731); 
 data3 <= my_rom(3086); 
 data4 <= my_rom(4441); 
 data5 <= my_rom(5796); 
 data6 <= my_rom(7151); 
 data7 <= my_rom(8506); 
 data8 <= my_rom(9861); 
 data9 <= my_rom(11216); 
 data10 <= my_rom(12571);
when "00101111001" => 
 data1 <= my_rom(377); 
 data2 <= my_rom(1732); 
 data3 <= my_rom(3087); 
 data4 <= my_rom(4442); 
 data5 <= my_rom(5797); 
 data6 <= my_rom(7152); 
 data7 <= my_rom(8507); 
 data8 <= my_rom(9862); 
 data9 <= my_rom(11217); 
 data10 <= my_rom(12572);
when "00101111010" => 
 data1 <= my_rom(378); 
 data2 <= my_rom(1733); 
 data3 <= my_rom(3088); 
 data4 <= my_rom(4443); 
 data5 <= my_rom(5798); 
 data6 <= my_rom(7153); 
 data7 <= my_rom(8508); 
 data8 <= my_rom(9863); 
 data9 <= my_rom(11218); 
 data10 <= my_rom(12573);
when "00101111011" => 
 data1 <= my_rom(379); 
 data2 <= my_rom(1734); 
 data3 <= my_rom(3089); 
 data4 <= my_rom(4444); 
 data5 <= my_rom(5799); 
 data6 <= my_rom(7154); 
 data7 <= my_rom(8509); 
 data8 <= my_rom(9864); 
 data9 <= my_rom(11219); 
 data10 <= my_rom(12574);
when "00101111100" => 
 data1 <= my_rom(380); 
 data2 <= my_rom(1735); 
 data3 <= my_rom(3090); 
 data4 <= my_rom(4445); 
 data5 <= my_rom(5800); 
 data6 <= my_rom(7155); 
 data7 <= my_rom(8510); 
 data8 <= my_rom(9865); 
 data9 <= my_rom(11220); 
 data10 <= my_rom(12575);
when "00101111101" => 
 data1 <= my_rom(381); 
 data2 <= my_rom(1736); 
 data3 <= my_rom(3091); 
 data4 <= my_rom(4446); 
 data5 <= my_rom(5801); 
 data6 <= my_rom(7156); 
 data7 <= my_rom(8511); 
 data8 <= my_rom(9866); 
 data9 <= my_rom(11221); 
 data10 <= my_rom(12576);
when "00101111110" => 
 data1 <= my_rom(382); 
 data2 <= my_rom(1737); 
 data3 <= my_rom(3092); 
 data4 <= my_rom(4447); 
 data5 <= my_rom(5802); 
 data6 <= my_rom(7157); 
 data7 <= my_rom(8512); 
 data8 <= my_rom(9867); 
 data9 <= my_rom(11222); 
 data10 <= my_rom(12577);
when "00101111111" => 
 data1 <= my_rom(383); 
 data2 <= my_rom(1738); 
 data3 <= my_rom(3093); 
 data4 <= my_rom(4448); 
 data5 <= my_rom(5803); 
 data6 <= my_rom(7158); 
 data7 <= my_rom(8513); 
 data8 <= my_rom(9868); 
 data9 <= my_rom(11223); 
 data10 <= my_rom(12578);
when "00110000000" => 
 data1 <= my_rom(384); 
 data2 <= my_rom(1739); 
 data3 <= my_rom(3094); 
 data4 <= my_rom(4449); 
 data5 <= my_rom(5804); 
 data6 <= my_rom(7159); 
 data7 <= my_rom(8514); 
 data8 <= my_rom(9869); 
 data9 <= my_rom(11224); 
 data10 <= my_rom(12579);
when "00110000001" => 
 data1 <= my_rom(385); 
 data2 <= my_rom(1740); 
 data3 <= my_rom(3095); 
 data4 <= my_rom(4450); 
 data5 <= my_rom(5805); 
 data6 <= my_rom(7160); 
 data7 <= my_rom(8515); 
 data8 <= my_rom(9870); 
 data9 <= my_rom(11225); 
 data10 <= my_rom(12580);
when "00110000010" => 
 data1 <= my_rom(386); 
 data2 <= my_rom(1741); 
 data3 <= my_rom(3096); 
 data4 <= my_rom(4451); 
 data5 <= my_rom(5806); 
 data6 <= my_rom(7161); 
 data7 <= my_rom(8516); 
 data8 <= my_rom(9871); 
 data9 <= my_rom(11226); 
 data10 <= my_rom(12581);
when "00110000011" => 
 data1 <= my_rom(387); 
 data2 <= my_rom(1742); 
 data3 <= my_rom(3097); 
 data4 <= my_rom(4452); 
 data5 <= my_rom(5807); 
 data6 <= my_rom(7162); 
 data7 <= my_rom(8517); 
 data8 <= my_rom(9872); 
 data9 <= my_rom(11227); 
 data10 <= my_rom(12582);
when "00110000100" => 
 data1 <= my_rom(388); 
 data2 <= my_rom(1743); 
 data3 <= my_rom(3098); 
 data4 <= my_rom(4453); 
 data5 <= my_rom(5808); 
 data6 <= my_rom(7163); 
 data7 <= my_rom(8518); 
 data8 <= my_rom(9873); 
 data9 <= my_rom(11228); 
 data10 <= my_rom(12583);
when "00110000101" => 
 data1 <= my_rom(389); 
 data2 <= my_rom(1744); 
 data3 <= my_rom(3099); 
 data4 <= my_rom(4454); 
 data5 <= my_rom(5809); 
 data6 <= my_rom(7164); 
 data7 <= my_rom(8519); 
 data8 <= my_rom(9874); 
 data9 <= my_rom(11229); 
 data10 <= my_rom(12584);
when "00110000110" => 
 data1 <= my_rom(390); 
 data2 <= my_rom(1745); 
 data3 <= my_rom(3100); 
 data4 <= my_rom(4455); 
 data5 <= my_rom(5810); 
 data6 <= my_rom(7165); 
 data7 <= my_rom(8520); 
 data8 <= my_rom(9875); 
 data9 <= my_rom(11230); 
 data10 <= my_rom(12585);
when "00110000111" => 
 data1 <= my_rom(391); 
 data2 <= my_rom(1746); 
 data3 <= my_rom(3101); 
 data4 <= my_rom(4456); 
 data5 <= my_rom(5811); 
 data6 <= my_rom(7166); 
 data7 <= my_rom(8521); 
 data8 <= my_rom(9876); 
 data9 <= my_rom(11231); 
 data10 <= my_rom(12586);
when "00110001000" => 
 data1 <= my_rom(392); 
 data2 <= my_rom(1747); 
 data3 <= my_rom(3102); 
 data4 <= my_rom(4457); 
 data5 <= my_rom(5812); 
 data6 <= my_rom(7167); 
 data7 <= my_rom(8522); 
 data8 <= my_rom(9877); 
 data9 <= my_rom(11232); 
 data10 <= my_rom(12587);
when "00110001001" => 
 data1 <= my_rom(393); 
 data2 <= my_rom(1748); 
 data3 <= my_rom(3103); 
 data4 <= my_rom(4458); 
 data5 <= my_rom(5813); 
 data6 <= my_rom(7168); 
 data7 <= my_rom(8523); 
 data8 <= my_rom(9878); 
 data9 <= my_rom(11233); 
 data10 <= my_rom(12588);
when "00110001010" => 
 data1 <= my_rom(394); 
 data2 <= my_rom(1749); 
 data3 <= my_rom(3104); 
 data4 <= my_rom(4459); 
 data5 <= my_rom(5814); 
 data6 <= my_rom(7169); 
 data7 <= my_rom(8524); 
 data8 <= my_rom(9879); 
 data9 <= my_rom(11234); 
 data10 <= my_rom(12589);
when "00110001011" => 
 data1 <= my_rom(395); 
 data2 <= my_rom(1750); 
 data3 <= my_rom(3105); 
 data4 <= my_rom(4460); 
 data5 <= my_rom(5815); 
 data6 <= my_rom(7170); 
 data7 <= my_rom(8525); 
 data8 <= my_rom(9880); 
 data9 <= my_rom(11235); 
 data10 <= my_rom(12590);
when "00110001100" => 
 data1 <= my_rom(396); 
 data2 <= my_rom(1751); 
 data3 <= my_rom(3106); 
 data4 <= my_rom(4461); 
 data5 <= my_rom(5816); 
 data6 <= my_rom(7171); 
 data7 <= my_rom(8526); 
 data8 <= my_rom(9881); 
 data9 <= my_rom(11236); 
 data10 <= my_rom(12591);
when "00110001101" => 
 data1 <= my_rom(397); 
 data2 <= my_rom(1752); 
 data3 <= my_rom(3107); 
 data4 <= my_rom(4462); 
 data5 <= my_rom(5817); 
 data6 <= my_rom(7172); 
 data7 <= my_rom(8527); 
 data8 <= my_rom(9882); 
 data9 <= my_rom(11237); 
 data10 <= my_rom(12592);
when "00110001110" => 
 data1 <= my_rom(398); 
 data2 <= my_rom(1753); 
 data3 <= my_rom(3108); 
 data4 <= my_rom(4463); 
 data5 <= my_rom(5818); 
 data6 <= my_rom(7173); 
 data7 <= my_rom(8528); 
 data8 <= my_rom(9883); 
 data9 <= my_rom(11238); 
 data10 <= my_rom(12593);
when "00110001111" => 
 data1 <= my_rom(399); 
 data2 <= my_rom(1754); 
 data3 <= my_rom(3109); 
 data4 <= my_rom(4464); 
 data5 <= my_rom(5819); 
 data6 <= my_rom(7174); 
 data7 <= my_rom(8529); 
 data8 <= my_rom(9884); 
 data9 <= my_rom(11239); 
 data10 <= my_rom(12594);
when "00110010000" => 
 data1 <= my_rom(400); 
 data2 <= my_rom(1755); 
 data3 <= my_rom(3110); 
 data4 <= my_rom(4465); 
 data5 <= my_rom(5820); 
 data6 <= my_rom(7175); 
 data7 <= my_rom(8530); 
 data8 <= my_rom(9885); 
 data9 <= my_rom(11240); 
 data10 <= my_rom(12595);
when "00110010001" => 
 data1 <= my_rom(401); 
 data2 <= my_rom(1756); 
 data3 <= my_rom(3111); 
 data4 <= my_rom(4466); 
 data5 <= my_rom(5821); 
 data6 <= my_rom(7176); 
 data7 <= my_rom(8531); 
 data8 <= my_rom(9886); 
 data9 <= my_rom(11241); 
 data10 <= my_rom(12596);
when "00110010010" => 
 data1 <= my_rom(402); 
 data2 <= my_rom(1757); 
 data3 <= my_rom(3112); 
 data4 <= my_rom(4467); 
 data5 <= my_rom(5822); 
 data6 <= my_rom(7177); 
 data7 <= my_rom(8532); 
 data8 <= my_rom(9887); 
 data9 <= my_rom(11242); 
 data10 <= my_rom(12597);
when "00110010011" => 
 data1 <= my_rom(403); 
 data2 <= my_rom(1758); 
 data3 <= my_rom(3113); 
 data4 <= my_rom(4468); 
 data5 <= my_rom(5823); 
 data6 <= my_rom(7178); 
 data7 <= my_rom(8533); 
 data8 <= my_rom(9888); 
 data9 <= my_rom(11243); 
 data10 <= my_rom(12598);
when "00110010100" => 
 data1 <= my_rom(404); 
 data2 <= my_rom(1759); 
 data3 <= my_rom(3114); 
 data4 <= my_rom(4469); 
 data5 <= my_rom(5824); 
 data6 <= my_rom(7179); 
 data7 <= my_rom(8534); 
 data8 <= my_rom(9889); 
 data9 <= my_rom(11244); 
 data10 <= my_rom(12599);
when "00110010101" => 
 data1 <= my_rom(405); 
 data2 <= my_rom(1760); 
 data3 <= my_rom(3115); 
 data4 <= my_rom(4470); 
 data5 <= my_rom(5825); 
 data6 <= my_rom(7180); 
 data7 <= my_rom(8535); 
 data8 <= my_rom(9890); 
 data9 <= my_rom(11245); 
 data10 <= my_rom(12600);
when "00110010110" => 
 data1 <= my_rom(406); 
 data2 <= my_rom(1761); 
 data3 <= my_rom(3116); 
 data4 <= my_rom(4471); 
 data5 <= my_rom(5826); 
 data6 <= my_rom(7181); 
 data7 <= my_rom(8536); 
 data8 <= my_rom(9891); 
 data9 <= my_rom(11246); 
 data10 <= my_rom(12601);
when "00110010111" => 
 data1 <= my_rom(407); 
 data2 <= my_rom(1762); 
 data3 <= my_rom(3117); 
 data4 <= my_rom(4472); 
 data5 <= my_rom(5827); 
 data6 <= my_rom(7182); 
 data7 <= my_rom(8537); 
 data8 <= my_rom(9892); 
 data9 <= my_rom(11247); 
 data10 <= my_rom(12602);
when "00110011000" => 
 data1 <= my_rom(408); 
 data2 <= my_rom(1763); 
 data3 <= my_rom(3118); 
 data4 <= my_rom(4473); 
 data5 <= my_rom(5828); 
 data6 <= my_rom(7183); 
 data7 <= my_rom(8538); 
 data8 <= my_rom(9893); 
 data9 <= my_rom(11248); 
 data10 <= my_rom(12603);
when "00110011001" => 
 data1 <= my_rom(409); 
 data2 <= my_rom(1764); 
 data3 <= my_rom(3119); 
 data4 <= my_rom(4474); 
 data5 <= my_rom(5829); 
 data6 <= my_rom(7184); 
 data7 <= my_rom(8539); 
 data8 <= my_rom(9894); 
 data9 <= my_rom(11249); 
 data10 <= my_rom(12604);
when "00110011010" => 
 data1 <= my_rom(410); 
 data2 <= my_rom(1765); 
 data3 <= my_rom(3120); 
 data4 <= my_rom(4475); 
 data5 <= my_rom(5830); 
 data6 <= my_rom(7185); 
 data7 <= my_rom(8540); 
 data8 <= my_rom(9895); 
 data9 <= my_rom(11250); 
 data10 <= my_rom(12605);
when "00110011011" => 
 data1 <= my_rom(411); 
 data2 <= my_rom(1766); 
 data3 <= my_rom(3121); 
 data4 <= my_rom(4476); 
 data5 <= my_rom(5831); 
 data6 <= my_rom(7186); 
 data7 <= my_rom(8541); 
 data8 <= my_rom(9896); 
 data9 <= my_rom(11251); 
 data10 <= my_rom(12606);
when "00110011100" => 
 data1 <= my_rom(412); 
 data2 <= my_rom(1767); 
 data3 <= my_rom(3122); 
 data4 <= my_rom(4477); 
 data5 <= my_rom(5832); 
 data6 <= my_rom(7187); 
 data7 <= my_rom(8542); 
 data8 <= my_rom(9897); 
 data9 <= my_rom(11252); 
 data10 <= my_rom(12607);
when "00110011101" => 
 data1 <= my_rom(413); 
 data2 <= my_rom(1768); 
 data3 <= my_rom(3123); 
 data4 <= my_rom(4478); 
 data5 <= my_rom(5833); 
 data6 <= my_rom(7188); 
 data7 <= my_rom(8543); 
 data8 <= my_rom(9898); 
 data9 <= my_rom(11253); 
 data10 <= my_rom(12608);
when "00110011110" => 
 data1 <= my_rom(414); 
 data2 <= my_rom(1769); 
 data3 <= my_rom(3124); 
 data4 <= my_rom(4479); 
 data5 <= my_rom(5834); 
 data6 <= my_rom(7189); 
 data7 <= my_rom(8544); 
 data8 <= my_rom(9899); 
 data9 <= my_rom(11254); 
 data10 <= my_rom(12609);
when "00110011111" => 
 data1 <= my_rom(415); 
 data2 <= my_rom(1770); 
 data3 <= my_rom(3125); 
 data4 <= my_rom(4480); 
 data5 <= my_rom(5835); 
 data6 <= my_rom(7190); 
 data7 <= my_rom(8545); 
 data8 <= my_rom(9900); 
 data9 <= my_rom(11255); 
 data10 <= my_rom(12610);
when "00110100000" => 
 data1 <= my_rom(416); 
 data2 <= my_rom(1771); 
 data3 <= my_rom(3126); 
 data4 <= my_rom(4481); 
 data5 <= my_rom(5836); 
 data6 <= my_rom(7191); 
 data7 <= my_rom(8546); 
 data8 <= my_rom(9901); 
 data9 <= my_rom(11256); 
 data10 <= my_rom(12611);
when "00110100001" => 
 data1 <= my_rom(417); 
 data2 <= my_rom(1772); 
 data3 <= my_rom(3127); 
 data4 <= my_rom(4482); 
 data5 <= my_rom(5837); 
 data6 <= my_rom(7192); 
 data7 <= my_rom(8547); 
 data8 <= my_rom(9902); 
 data9 <= my_rom(11257); 
 data10 <= my_rom(12612);
when "00110100010" => 
 data1 <= my_rom(418); 
 data2 <= my_rom(1773); 
 data3 <= my_rom(3128); 
 data4 <= my_rom(4483); 
 data5 <= my_rom(5838); 
 data6 <= my_rom(7193); 
 data7 <= my_rom(8548); 
 data8 <= my_rom(9903); 
 data9 <= my_rom(11258); 
 data10 <= my_rom(12613);
when "00110100011" => 
 data1 <= my_rom(419); 
 data2 <= my_rom(1774); 
 data3 <= my_rom(3129); 
 data4 <= my_rom(4484); 
 data5 <= my_rom(5839); 
 data6 <= my_rom(7194); 
 data7 <= my_rom(8549); 
 data8 <= my_rom(9904); 
 data9 <= my_rom(11259); 
 data10 <= my_rom(12614);
when "00110100100" => 
 data1 <= my_rom(420); 
 data2 <= my_rom(1775); 
 data3 <= my_rom(3130); 
 data4 <= my_rom(4485); 
 data5 <= my_rom(5840); 
 data6 <= my_rom(7195); 
 data7 <= my_rom(8550); 
 data8 <= my_rom(9905); 
 data9 <= my_rom(11260); 
 data10 <= my_rom(12615);
when "00110100101" => 
 data1 <= my_rom(421); 
 data2 <= my_rom(1776); 
 data3 <= my_rom(3131); 
 data4 <= my_rom(4486); 
 data5 <= my_rom(5841); 
 data6 <= my_rom(7196); 
 data7 <= my_rom(8551); 
 data8 <= my_rom(9906); 
 data9 <= my_rom(11261); 
 data10 <= my_rom(12616);
when "00110100110" => 
 data1 <= my_rom(422); 
 data2 <= my_rom(1777); 
 data3 <= my_rom(3132); 
 data4 <= my_rom(4487); 
 data5 <= my_rom(5842); 
 data6 <= my_rom(7197); 
 data7 <= my_rom(8552); 
 data8 <= my_rom(9907); 
 data9 <= my_rom(11262); 
 data10 <= my_rom(12617);
when "00110100111" => 
 data1 <= my_rom(423); 
 data2 <= my_rom(1778); 
 data3 <= my_rom(3133); 
 data4 <= my_rom(4488); 
 data5 <= my_rom(5843); 
 data6 <= my_rom(7198); 
 data7 <= my_rom(8553); 
 data8 <= my_rom(9908); 
 data9 <= my_rom(11263); 
 data10 <= my_rom(12618);
when "00110101000" => 
 data1 <= my_rom(424); 
 data2 <= my_rom(1779); 
 data3 <= my_rom(3134); 
 data4 <= my_rom(4489); 
 data5 <= my_rom(5844); 
 data6 <= my_rom(7199); 
 data7 <= my_rom(8554); 
 data8 <= my_rom(9909); 
 data9 <= my_rom(11264); 
 data10 <= my_rom(12619);
when "00110101001" => 
 data1 <= my_rom(425); 
 data2 <= my_rom(1780); 
 data3 <= my_rom(3135); 
 data4 <= my_rom(4490); 
 data5 <= my_rom(5845); 
 data6 <= my_rom(7200); 
 data7 <= my_rom(8555); 
 data8 <= my_rom(9910); 
 data9 <= my_rom(11265); 
 data10 <= my_rom(12620);
when "00110101010" => 
 data1 <= my_rom(426); 
 data2 <= my_rom(1781); 
 data3 <= my_rom(3136); 
 data4 <= my_rom(4491); 
 data5 <= my_rom(5846); 
 data6 <= my_rom(7201); 
 data7 <= my_rom(8556); 
 data8 <= my_rom(9911); 
 data9 <= my_rom(11266); 
 data10 <= my_rom(12621);
when "00110101011" => 
 data1 <= my_rom(427); 
 data2 <= my_rom(1782); 
 data3 <= my_rom(3137); 
 data4 <= my_rom(4492); 
 data5 <= my_rom(5847); 
 data6 <= my_rom(7202); 
 data7 <= my_rom(8557); 
 data8 <= my_rom(9912); 
 data9 <= my_rom(11267); 
 data10 <= my_rom(12622);
when "00110101100" => 
 data1 <= my_rom(428); 
 data2 <= my_rom(1783); 
 data3 <= my_rom(3138); 
 data4 <= my_rom(4493); 
 data5 <= my_rom(5848); 
 data6 <= my_rom(7203); 
 data7 <= my_rom(8558); 
 data8 <= my_rom(9913); 
 data9 <= my_rom(11268); 
 data10 <= my_rom(12623);
when "00110101101" => 
 data1 <= my_rom(429); 
 data2 <= my_rom(1784); 
 data3 <= my_rom(3139); 
 data4 <= my_rom(4494); 
 data5 <= my_rom(5849); 
 data6 <= my_rom(7204); 
 data7 <= my_rom(8559); 
 data8 <= my_rom(9914); 
 data9 <= my_rom(11269); 
 data10 <= my_rom(12624);
when "00110101110" => 
 data1 <= my_rom(430); 
 data2 <= my_rom(1785); 
 data3 <= my_rom(3140); 
 data4 <= my_rom(4495); 
 data5 <= my_rom(5850); 
 data6 <= my_rom(7205); 
 data7 <= my_rom(8560); 
 data8 <= my_rom(9915); 
 data9 <= my_rom(11270); 
 data10 <= my_rom(12625);
when "00110101111" => 
 data1 <= my_rom(431); 
 data2 <= my_rom(1786); 
 data3 <= my_rom(3141); 
 data4 <= my_rom(4496); 
 data5 <= my_rom(5851); 
 data6 <= my_rom(7206); 
 data7 <= my_rom(8561); 
 data8 <= my_rom(9916); 
 data9 <= my_rom(11271); 
 data10 <= my_rom(12626);
when "00110110000" => 
 data1 <= my_rom(432); 
 data2 <= my_rom(1787); 
 data3 <= my_rom(3142); 
 data4 <= my_rom(4497); 
 data5 <= my_rom(5852); 
 data6 <= my_rom(7207); 
 data7 <= my_rom(8562); 
 data8 <= my_rom(9917); 
 data9 <= my_rom(11272); 
 data10 <= my_rom(12627);
when "00110110001" => 
 data1 <= my_rom(433); 
 data2 <= my_rom(1788); 
 data3 <= my_rom(3143); 
 data4 <= my_rom(4498); 
 data5 <= my_rom(5853); 
 data6 <= my_rom(7208); 
 data7 <= my_rom(8563); 
 data8 <= my_rom(9918); 
 data9 <= my_rom(11273); 
 data10 <= my_rom(12628);
when "00110110010" => 
 data1 <= my_rom(434); 
 data2 <= my_rom(1789); 
 data3 <= my_rom(3144); 
 data4 <= my_rom(4499); 
 data5 <= my_rom(5854); 
 data6 <= my_rom(7209); 
 data7 <= my_rom(8564); 
 data8 <= my_rom(9919); 
 data9 <= my_rom(11274); 
 data10 <= my_rom(12629);
when "00110110011" => 
 data1 <= my_rom(435); 
 data2 <= my_rom(1790); 
 data3 <= my_rom(3145); 
 data4 <= my_rom(4500); 
 data5 <= my_rom(5855); 
 data6 <= my_rom(7210); 
 data7 <= my_rom(8565); 
 data8 <= my_rom(9920); 
 data9 <= my_rom(11275); 
 data10 <= my_rom(12630);
when "00110110100" => 
 data1 <= my_rom(436); 
 data2 <= my_rom(1791); 
 data3 <= my_rom(3146); 
 data4 <= my_rom(4501); 
 data5 <= my_rom(5856); 
 data6 <= my_rom(7211); 
 data7 <= my_rom(8566); 
 data8 <= my_rom(9921); 
 data9 <= my_rom(11276); 
 data10 <= my_rom(12631);
when "00110110101" => 
 data1 <= my_rom(437); 
 data2 <= my_rom(1792); 
 data3 <= my_rom(3147); 
 data4 <= my_rom(4502); 
 data5 <= my_rom(5857); 
 data6 <= my_rom(7212); 
 data7 <= my_rom(8567); 
 data8 <= my_rom(9922); 
 data9 <= my_rom(11277); 
 data10 <= my_rom(12632);
when "00110110110" => 
 data1 <= my_rom(438); 
 data2 <= my_rom(1793); 
 data3 <= my_rom(3148); 
 data4 <= my_rom(4503); 
 data5 <= my_rom(5858); 
 data6 <= my_rom(7213); 
 data7 <= my_rom(8568); 
 data8 <= my_rom(9923); 
 data9 <= my_rom(11278); 
 data10 <= my_rom(12633);
when "00110110111" => 
 data1 <= my_rom(439); 
 data2 <= my_rom(1794); 
 data3 <= my_rom(3149); 
 data4 <= my_rom(4504); 
 data5 <= my_rom(5859); 
 data6 <= my_rom(7214); 
 data7 <= my_rom(8569); 
 data8 <= my_rom(9924); 
 data9 <= my_rom(11279); 
 data10 <= my_rom(12634);
when "00110111000" => 
 data1 <= my_rom(440); 
 data2 <= my_rom(1795); 
 data3 <= my_rom(3150); 
 data4 <= my_rom(4505); 
 data5 <= my_rom(5860); 
 data6 <= my_rom(7215); 
 data7 <= my_rom(8570); 
 data8 <= my_rom(9925); 
 data9 <= my_rom(11280); 
 data10 <= my_rom(12635);
when "00110111001" => 
 data1 <= my_rom(441); 
 data2 <= my_rom(1796); 
 data3 <= my_rom(3151); 
 data4 <= my_rom(4506); 
 data5 <= my_rom(5861); 
 data6 <= my_rom(7216); 
 data7 <= my_rom(8571); 
 data8 <= my_rom(9926); 
 data9 <= my_rom(11281); 
 data10 <= my_rom(12636);
when "00110111010" => 
 data1 <= my_rom(442); 
 data2 <= my_rom(1797); 
 data3 <= my_rom(3152); 
 data4 <= my_rom(4507); 
 data5 <= my_rom(5862); 
 data6 <= my_rom(7217); 
 data7 <= my_rom(8572); 
 data8 <= my_rom(9927); 
 data9 <= my_rom(11282); 
 data10 <= my_rom(12637);
when "00110111011" => 
 data1 <= my_rom(443); 
 data2 <= my_rom(1798); 
 data3 <= my_rom(3153); 
 data4 <= my_rom(4508); 
 data5 <= my_rom(5863); 
 data6 <= my_rom(7218); 
 data7 <= my_rom(8573); 
 data8 <= my_rom(9928); 
 data9 <= my_rom(11283); 
 data10 <= my_rom(12638);
when "00110111100" => 
 data1 <= my_rom(444); 
 data2 <= my_rom(1799); 
 data3 <= my_rom(3154); 
 data4 <= my_rom(4509); 
 data5 <= my_rom(5864); 
 data6 <= my_rom(7219); 
 data7 <= my_rom(8574); 
 data8 <= my_rom(9929); 
 data9 <= my_rom(11284); 
 data10 <= my_rom(12639);
when "00110111101" => 
 data1 <= my_rom(445); 
 data2 <= my_rom(1800); 
 data3 <= my_rom(3155); 
 data4 <= my_rom(4510); 
 data5 <= my_rom(5865); 
 data6 <= my_rom(7220); 
 data7 <= my_rom(8575); 
 data8 <= my_rom(9930); 
 data9 <= my_rom(11285); 
 data10 <= my_rom(12640);
when "00110111110" => 
 data1 <= my_rom(446); 
 data2 <= my_rom(1801); 
 data3 <= my_rom(3156); 
 data4 <= my_rom(4511); 
 data5 <= my_rom(5866); 
 data6 <= my_rom(7221); 
 data7 <= my_rom(8576); 
 data8 <= my_rom(9931); 
 data9 <= my_rom(11286); 
 data10 <= my_rom(12641);
when "00110111111" => 
 data1 <= my_rom(447); 
 data2 <= my_rom(1802); 
 data3 <= my_rom(3157); 
 data4 <= my_rom(4512); 
 data5 <= my_rom(5867); 
 data6 <= my_rom(7222); 
 data7 <= my_rom(8577); 
 data8 <= my_rom(9932); 
 data9 <= my_rom(11287); 
 data10 <= my_rom(12642);
when "00111000000" => 
 data1 <= my_rom(448); 
 data2 <= my_rom(1803); 
 data3 <= my_rom(3158); 
 data4 <= my_rom(4513); 
 data5 <= my_rom(5868); 
 data6 <= my_rom(7223); 
 data7 <= my_rom(8578); 
 data8 <= my_rom(9933); 
 data9 <= my_rom(11288); 
 data10 <= my_rom(12643);
when "00111000001" => 
 data1 <= my_rom(449); 
 data2 <= my_rom(1804); 
 data3 <= my_rom(3159); 
 data4 <= my_rom(4514); 
 data5 <= my_rom(5869); 
 data6 <= my_rom(7224); 
 data7 <= my_rom(8579); 
 data8 <= my_rom(9934); 
 data9 <= my_rom(11289); 
 data10 <= my_rom(12644);
when "00111000010" => 
 data1 <= my_rom(450); 
 data2 <= my_rom(1805); 
 data3 <= my_rom(3160); 
 data4 <= my_rom(4515); 
 data5 <= my_rom(5870); 
 data6 <= my_rom(7225); 
 data7 <= my_rom(8580); 
 data8 <= my_rom(9935); 
 data9 <= my_rom(11290); 
 data10 <= my_rom(12645);
when "00111000011" => 
 data1 <= my_rom(451); 
 data2 <= my_rom(1806); 
 data3 <= my_rom(3161); 
 data4 <= my_rom(4516); 
 data5 <= my_rom(5871); 
 data6 <= my_rom(7226); 
 data7 <= my_rom(8581); 
 data8 <= my_rom(9936); 
 data9 <= my_rom(11291); 
 data10 <= my_rom(12646);
when "00111000100" => 
 data1 <= my_rom(452); 
 data2 <= my_rom(1807); 
 data3 <= my_rom(3162); 
 data4 <= my_rom(4517); 
 data5 <= my_rom(5872); 
 data6 <= my_rom(7227); 
 data7 <= my_rom(8582); 
 data8 <= my_rom(9937); 
 data9 <= my_rom(11292); 
 data10 <= my_rom(12647);
when "00111000101" => 
 data1 <= my_rom(453); 
 data2 <= my_rom(1808); 
 data3 <= my_rom(3163); 
 data4 <= my_rom(4518); 
 data5 <= my_rom(5873); 
 data6 <= my_rom(7228); 
 data7 <= my_rom(8583); 
 data8 <= my_rom(9938); 
 data9 <= my_rom(11293); 
 data10 <= my_rom(12648);
when "00111000110" => 
 data1 <= my_rom(454); 
 data2 <= my_rom(1809); 
 data3 <= my_rom(3164); 
 data4 <= my_rom(4519); 
 data5 <= my_rom(5874); 
 data6 <= my_rom(7229); 
 data7 <= my_rom(8584); 
 data8 <= my_rom(9939); 
 data9 <= my_rom(11294); 
 data10 <= my_rom(12649);
when "00111000111" => 
 data1 <= my_rom(455); 
 data2 <= my_rom(1810); 
 data3 <= my_rom(3165); 
 data4 <= my_rom(4520); 
 data5 <= my_rom(5875); 
 data6 <= my_rom(7230); 
 data7 <= my_rom(8585); 
 data8 <= my_rom(9940); 
 data9 <= my_rom(11295); 
 data10 <= my_rom(12650);
when "00111001000" => 
 data1 <= my_rom(456); 
 data2 <= my_rom(1811); 
 data3 <= my_rom(3166); 
 data4 <= my_rom(4521); 
 data5 <= my_rom(5876); 
 data6 <= my_rom(7231); 
 data7 <= my_rom(8586); 
 data8 <= my_rom(9941); 
 data9 <= my_rom(11296); 
 data10 <= my_rom(12651);
when "00111001001" => 
 data1 <= my_rom(457); 
 data2 <= my_rom(1812); 
 data3 <= my_rom(3167); 
 data4 <= my_rom(4522); 
 data5 <= my_rom(5877); 
 data6 <= my_rom(7232); 
 data7 <= my_rom(8587); 
 data8 <= my_rom(9942); 
 data9 <= my_rom(11297); 
 data10 <= my_rom(12652);
when "00111001010" => 
 data1 <= my_rom(458); 
 data2 <= my_rom(1813); 
 data3 <= my_rom(3168); 
 data4 <= my_rom(4523); 
 data5 <= my_rom(5878); 
 data6 <= my_rom(7233); 
 data7 <= my_rom(8588); 
 data8 <= my_rom(9943); 
 data9 <= my_rom(11298); 
 data10 <= my_rom(12653);
when "00111001011" => 
 data1 <= my_rom(459); 
 data2 <= my_rom(1814); 
 data3 <= my_rom(3169); 
 data4 <= my_rom(4524); 
 data5 <= my_rom(5879); 
 data6 <= my_rom(7234); 
 data7 <= my_rom(8589); 
 data8 <= my_rom(9944); 
 data9 <= my_rom(11299); 
 data10 <= my_rom(12654);
when "00111001100" => 
 data1 <= my_rom(460); 
 data2 <= my_rom(1815); 
 data3 <= my_rom(3170); 
 data4 <= my_rom(4525); 
 data5 <= my_rom(5880); 
 data6 <= my_rom(7235); 
 data7 <= my_rom(8590); 
 data8 <= my_rom(9945); 
 data9 <= my_rom(11300); 
 data10 <= my_rom(12655);
when "00111001101" => 
 data1 <= my_rom(461); 
 data2 <= my_rom(1816); 
 data3 <= my_rom(3171); 
 data4 <= my_rom(4526); 
 data5 <= my_rom(5881); 
 data6 <= my_rom(7236); 
 data7 <= my_rom(8591); 
 data8 <= my_rom(9946); 
 data9 <= my_rom(11301); 
 data10 <= my_rom(12656);
when "00111001110" => 
 data1 <= my_rom(462); 
 data2 <= my_rom(1817); 
 data3 <= my_rom(3172); 
 data4 <= my_rom(4527); 
 data5 <= my_rom(5882); 
 data6 <= my_rom(7237); 
 data7 <= my_rom(8592); 
 data8 <= my_rom(9947); 
 data9 <= my_rom(11302); 
 data10 <= my_rom(12657);
when "00111001111" => 
 data1 <= my_rom(463); 
 data2 <= my_rom(1818); 
 data3 <= my_rom(3173); 
 data4 <= my_rom(4528); 
 data5 <= my_rom(5883); 
 data6 <= my_rom(7238); 
 data7 <= my_rom(8593); 
 data8 <= my_rom(9948); 
 data9 <= my_rom(11303); 
 data10 <= my_rom(12658);
when "00111010000" => 
 data1 <= my_rom(464); 
 data2 <= my_rom(1819); 
 data3 <= my_rom(3174); 
 data4 <= my_rom(4529); 
 data5 <= my_rom(5884); 
 data6 <= my_rom(7239); 
 data7 <= my_rom(8594); 
 data8 <= my_rom(9949); 
 data9 <= my_rom(11304); 
 data10 <= my_rom(12659);
when "00111010001" => 
 data1 <= my_rom(465); 
 data2 <= my_rom(1820); 
 data3 <= my_rom(3175); 
 data4 <= my_rom(4530); 
 data5 <= my_rom(5885); 
 data6 <= my_rom(7240); 
 data7 <= my_rom(8595); 
 data8 <= my_rom(9950); 
 data9 <= my_rom(11305); 
 data10 <= my_rom(12660);
when "00111010010" => 
 data1 <= my_rom(466); 
 data2 <= my_rom(1821); 
 data3 <= my_rom(3176); 
 data4 <= my_rom(4531); 
 data5 <= my_rom(5886); 
 data6 <= my_rom(7241); 
 data7 <= my_rom(8596); 
 data8 <= my_rom(9951); 
 data9 <= my_rom(11306); 
 data10 <= my_rom(12661);
when "00111010011" => 
 data1 <= my_rom(467); 
 data2 <= my_rom(1822); 
 data3 <= my_rom(3177); 
 data4 <= my_rom(4532); 
 data5 <= my_rom(5887); 
 data6 <= my_rom(7242); 
 data7 <= my_rom(8597); 
 data8 <= my_rom(9952); 
 data9 <= my_rom(11307); 
 data10 <= my_rom(12662);
when "00111010100" => 
 data1 <= my_rom(468); 
 data2 <= my_rom(1823); 
 data3 <= my_rom(3178); 
 data4 <= my_rom(4533); 
 data5 <= my_rom(5888); 
 data6 <= my_rom(7243); 
 data7 <= my_rom(8598); 
 data8 <= my_rom(9953); 
 data9 <= my_rom(11308); 
 data10 <= my_rom(12663);
when "00111010101" => 
 data1 <= my_rom(469); 
 data2 <= my_rom(1824); 
 data3 <= my_rom(3179); 
 data4 <= my_rom(4534); 
 data5 <= my_rom(5889); 
 data6 <= my_rom(7244); 
 data7 <= my_rom(8599); 
 data8 <= my_rom(9954); 
 data9 <= my_rom(11309); 
 data10 <= my_rom(12664);
when "00111010110" => 
 data1 <= my_rom(470); 
 data2 <= my_rom(1825); 
 data3 <= my_rom(3180); 
 data4 <= my_rom(4535); 
 data5 <= my_rom(5890); 
 data6 <= my_rom(7245); 
 data7 <= my_rom(8600); 
 data8 <= my_rom(9955); 
 data9 <= my_rom(11310); 
 data10 <= my_rom(12665);
when "00111010111" => 
 data1 <= my_rom(471); 
 data2 <= my_rom(1826); 
 data3 <= my_rom(3181); 
 data4 <= my_rom(4536); 
 data5 <= my_rom(5891); 
 data6 <= my_rom(7246); 
 data7 <= my_rom(8601); 
 data8 <= my_rom(9956); 
 data9 <= my_rom(11311); 
 data10 <= my_rom(12666);
when "00111011000" => 
 data1 <= my_rom(472); 
 data2 <= my_rom(1827); 
 data3 <= my_rom(3182); 
 data4 <= my_rom(4537); 
 data5 <= my_rom(5892); 
 data6 <= my_rom(7247); 
 data7 <= my_rom(8602); 
 data8 <= my_rom(9957); 
 data9 <= my_rom(11312); 
 data10 <= my_rom(12667);
when "00111011001" => 
 data1 <= my_rom(473); 
 data2 <= my_rom(1828); 
 data3 <= my_rom(3183); 
 data4 <= my_rom(4538); 
 data5 <= my_rom(5893); 
 data6 <= my_rom(7248); 
 data7 <= my_rom(8603); 
 data8 <= my_rom(9958); 
 data9 <= my_rom(11313); 
 data10 <= my_rom(12668);
when "00111011010" => 
 data1 <= my_rom(474); 
 data2 <= my_rom(1829); 
 data3 <= my_rom(3184); 
 data4 <= my_rom(4539); 
 data5 <= my_rom(5894); 
 data6 <= my_rom(7249); 
 data7 <= my_rom(8604); 
 data8 <= my_rom(9959); 
 data9 <= my_rom(11314); 
 data10 <= my_rom(12669);
when "00111011011" => 
 data1 <= my_rom(475); 
 data2 <= my_rom(1830); 
 data3 <= my_rom(3185); 
 data4 <= my_rom(4540); 
 data5 <= my_rom(5895); 
 data6 <= my_rom(7250); 
 data7 <= my_rom(8605); 
 data8 <= my_rom(9960); 
 data9 <= my_rom(11315); 
 data10 <= my_rom(12670);
when "00111011100" => 
 data1 <= my_rom(476); 
 data2 <= my_rom(1831); 
 data3 <= my_rom(3186); 
 data4 <= my_rom(4541); 
 data5 <= my_rom(5896); 
 data6 <= my_rom(7251); 
 data7 <= my_rom(8606); 
 data8 <= my_rom(9961); 
 data9 <= my_rom(11316); 
 data10 <= my_rom(12671);
when "00111011101" => 
 data1 <= my_rom(477); 
 data2 <= my_rom(1832); 
 data3 <= my_rom(3187); 
 data4 <= my_rom(4542); 
 data5 <= my_rom(5897); 
 data6 <= my_rom(7252); 
 data7 <= my_rom(8607); 
 data8 <= my_rom(9962); 
 data9 <= my_rom(11317); 
 data10 <= my_rom(12672);
when "00111011110" => 
 data1 <= my_rom(478); 
 data2 <= my_rom(1833); 
 data3 <= my_rom(3188); 
 data4 <= my_rom(4543); 
 data5 <= my_rom(5898); 
 data6 <= my_rom(7253); 
 data7 <= my_rom(8608); 
 data8 <= my_rom(9963); 
 data9 <= my_rom(11318); 
 data10 <= my_rom(12673);
when "00111011111" => 
 data1 <= my_rom(479); 
 data2 <= my_rom(1834); 
 data3 <= my_rom(3189); 
 data4 <= my_rom(4544); 
 data5 <= my_rom(5899); 
 data6 <= my_rom(7254); 
 data7 <= my_rom(8609); 
 data8 <= my_rom(9964); 
 data9 <= my_rom(11319); 
 data10 <= my_rom(12674);
when "00111100000" => 
 data1 <= my_rom(480); 
 data2 <= my_rom(1835); 
 data3 <= my_rom(3190); 
 data4 <= my_rom(4545); 
 data5 <= my_rom(5900); 
 data6 <= my_rom(7255); 
 data7 <= my_rom(8610); 
 data8 <= my_rom(9965); 
 data9 <= my_rom(11320); 
 data10 <= my_rom(12675);
when "00111100001" => 
 data1 <= my_rom(481); 
 data2 <= my_rom(1836); 
 data3 <= my_rom(3191); 
 data4 <= my_rom(4546); 
 data5 <= my_rom(5901); 
 data6 <= my_rom(7256); 
 data7 <= my_rom(8611); 
 data8 <= my_rom(9966); 
 data9 <= my_rom(11321); 
 data10 <= my_rom(12676);
when "00111100010" => 
 data1 <= my_rom(482); 
 data2 <= my_rom(1837); 
 data3 <= my_rom(3192); 
 data4 <= my_rom(4547); 
 data5 <= my_rom(5902); 
 data6 <= my_rom(7257); 
 data7 <= my_rom(8612); 
 data8 <= my_rom(9967); 
 data9 <= my_rom(11322); 
 data10 <= my_rom(12677);
when "00111100011" => 
 data1 <= my_rom(483); 
 data2 <= my_rom(1838); 
 data3 <= my_rom(3193); 
 data4 <= my_rom(4548); 
 data5 <= my_rom(5903); 
 data6 <= my_rom(7258); 
 data7 <= my_rom(8613); 
 data8 <= my_rom(9968); 
 data9 <= my_rom(11323); 
 data10 <= my_rom(12678);
when "00111100100" => 
 data1 <= my_rom(484); 
 data2 <= my_rom(1839); 
 data3 <= my_rom(3194); 
 data4 <= my_rom(4549); 
 data5 <= my_rom(5904); 
 data6 <= my_rom(7259); 
 data7 <= my_rom(8614); 
 data8 <= my_rom(9969); 
 data9 <= my_rom(11324); 
 data10 <= my_rom(12679);
when "00111100101" => 
 data1 <= my_rom(485); 
 data2 <= my_rom(1840); 
 data3 <= my_rom(3195); 
 data4 <= my_rom(4550); 
 data5 <= my_rom(5905); 
 data6 <= my_rom(7260); 
 data7 <= my_rom(8615); 
 data8 <= my_rom(9970); 
 data9 <= my_rom(11325); 
 data10 <= my_rom(12680);
when "00111100110" => 
 data1 <= my_rom(486); 
 data2 <= my_rom(1841); 
 data3 <= my_rom(3196); 
 data4 <= my_rom(4551); 
 data5 <= my_rom(5906); 
 data6 <= my_rom(7261); 
 data7 <= my_rom(8616); 
 data8 <= my_rom(9971); 
 data9 <= my_rom(11326); 
 data10 <= my_rom(12681);
when "00111100111" => 
 data1 <= my_rom(487); 
 data2 <= my_rom(1842); 
 data3 <= my_rom(3197); 
 data4 <= my_rom(4552); 
 data5 <= my_rom(5907); 
 data6 <= my_rom(7262); 
 data7 <= my_rom(8617); 
 data8 <= my_rom(9972); 
 data9 <= my_rom(11327); 
 data10 <= my_rom(12682);
when "00111101000" => 
 data1 <= my_rom(488); 
 data2 <= my_rom(1843); 
 data3 <= my_rom(3198); 
 data4 <= my_rom(4553); 
 data5 <= my_rom(5908); 
 data6 <= my_rom(7263); 
 data7 <= my_rom(8618); 
 data8 <= my_rom(9973); 
 data9 <= my_rom(11328); 
 data10 <= my_rom(12683);
when "00111101001" => 
 data1 <= my_rom(489); 
 data2 <= my_rom(1844); 
 data3 <= my_rom(3199); 
 data4 <= my_rom(4554); 
 data5 <= my_rom(5909); 
 data6 <= my_rom(7264); 
 data7 <= my_rom(8619); 
 data8 <= my_rom(9974); 
 data9 <= my_rom(11329); 
 data10 <= my_rom(12684);
when "00111101010" => 
 data1 <= my_rom(490); 
 data2 <= my_rom(1845); 
 data3 <= my_rom(3200); 
 data4 <= my_rom(4555); 
 data5 <= my_rom(5910); 
 data6 <= my_rom(7265); 
 data7 <= my_rom(8620); 
 data8 <= my_rom(9975); 
 data9 <= my_rom(11330); 
 data10 <= my_rom(12685);
when "00111101011" => 
 data1 <= my_rom(491); 
 data2 <= my_rom(1846); 
 data3 <= my_rom(3201); 
 data4 <= my_rom(4556); 
 data5 <= my_rom(5911); 
 data6 <= my_rom(7266); 
 data7 <= my_rom(8621); 
 data8 <= my_rom(9976); 
 data9 <= my_rom(11331); 
 data10 <= my_rom(12686);
when "00111101100" => 
 data1 <= my_rom(492); 
 data2 <= my_rom(1847); 
 data3 <= my_rom(3202); 
 data4 <= my_rom(4557); 
 data5 <= my_rom(5912); 
 data6 <= my_rom(7267); 
 data7 <= my_rom(8622); 
 data8 <= my_rom(9977); 
 data9 <= my_rom(11332); 
 data10 <= my_rom(12687);
when "00111101101" => 
 data1 <= my_rom(493); 
 data2 <= my_rom(1848); 
 data3 <= my_rom(3203); 
 data4 <= my_rom(4558); 
 data5 <= my_rom(5913); 
 data6 <= my_rom(7268); 
 data7 <= my_rom(8623); 
 data8 <= my_rom(9978); 
 data9 <= my_rom(11333); 
 data10 <= my_rom(12688);
when "00111101110" => 
 data1 <= my_rom(494); 
 data2 <= my_rom(1849); 
 data3 <= my_rom(3204); 
 data4 <= my_rom(4559); 
 data5 <= my_rom(5914); 
 data6 <= my_rom(7269); 
 data7 <= my_rom(8624); 
 data8 <= my_rom(9979); 
 data9 <= my_rom(11334); 
 data10 <= my_rom(12689);
when "00111101111" => 
 data1 <= my_rom(495); 
 data2 <= my_rom(1850); 
 data3 <= my_rom(3205); 
 data4 <= my_rom(4560); 
 data5 <= my_rom(5915); 
 data6 <= my_rom(7270); 
 data7 <= my_rom(8625); 
 data8 <= my_rom(9980); 
 data9 <= my_rom(11335); 
 data10 <= my_rom(12690);
when "00111110000" => 
 data1 <= my_rom(496); 
 data2 <= my_rom(1851); 
 data3 <= my_rom(3206); 
 data4 <= my_rom(4561); 
 data5 <= my_rom(5916); 
 data6 <= my_rom(7271); 
 data7 <= my_rom(8626); 
 data8 <= my_rom(9981); 
 data9 <= my_rom(11336); 
 data10 <= my_rom(12691);
when "00111110001" => 
 data1 <= my_rom(497); 
 data2 <= my_rom(1852); 
 data3 <= my_rom(3207); 
 data4 <= my_rom(4562); 
 data5 <= my_rom(5917); 
 data6 <= my_rom(7272); 
 data7 <= my_rom(8627); 
 data8 <= my_rom(9982); 
 data9 <= my_rom(11337); 
 data10 <= my_rom(12692);
when "00111110010" => 
 data1 <= my_rom(498); 
 data2 <= my_rom(1853); 
 data3 <= my_rom(3208); 
 data4 <= my_rom(4563); 
 data5 <= my_rom(5918); 
 data6 <= my_rom(7273); 
 data7 <= my_rom(8628); 
 data8 <= my_rom(9983); 
 data9 <= my_rom(11338); 
 data10 <= my_rom(12693);
when "00111110011" => 
 data1 <= my_rom(499); 
 data2 <= my_rom(1854); 
 data3 <= my_rom(3209); 
 data4 <= my_rom(4564); 
 data5 <= my_rom(5919); 
 data6 <= my_rom(7274); 
 data7 <= my_rom(8629); 
 data8 <= my_rom(9984); 
 data9 <= my_rom(11339); 
 data10 <= my_rom(12694);
when "00111110100" => 
 data1 <= my_rom(500); 
 data2 <= my_rom(1855); 
 data3 <= my_rom(3210); 
 data4 <= my_rom(4565); 
 data5 <= my_rom(5920); 
 data6 <= my_rom(7275); 
 data7 <= my_rom(8630); 
 data8 <= my_rom(9985); 
 data9 <= my_rom(11340); 
 data10 <= my_rom(12695);
when "00111110101" => 
 data1 <= my_rom(501); 
 data2 <= my_rom(1856); 
 data3 <= my_rom(3211); 
 data4 <= my_rom(4566); 
 data5 <= my_rom(5921); 
 data6 <= my_rom(7276); 
 data7 <= my_rom(8631); 
 data8 <= my_rom(9986); 
 data9 <= my_rom(11341); 
 data10 <= my_rom(12696);
when "00111110110" => 
 data1 <= my_rom(502); 
 data2 <= my_rom(1857); 
 data3 <= my_rom(3212); 
 data4 <= my_rom(4567); 
 data5 <= my_rom(5922); 
 data6 <= my_rom(7277); 
 data7 <= my_rom(8632); 
 data8 <= my_rom(9987); 
 data9 <= my_rom(11342); 
 data10 <= my_rom(12697);
when "00111110111" => 
 data1 <= my_rom(503); 
 data2 <= my_rom(1858); 
 data3 <= my_rom(3213); 
 data4 <= my_rom(4568); 
 data5 <= my_rom(5923); 
 data6 <= my_rom(7278); 
 data7 <= my_rom(8633); 
 data8 <= my_rom(9988); 
 data9 <= my_rom(11343); 
 data10 <= my_rom(12698);
when "00111111000" => 
 data1 <= my_rom(504); 
 data2 <= my_rom(1859); 
 data3 <= my_rom(3214); 
 data4 <= my_rom(4569); 
 data5 <= my_rom(5924); 
 data6 <= my_rom(7279); 
 data7 <= my_rom(8634); 
 data8 <= my_rom(9989); 
 data9 <= my_rom(11344); 
 data10 <= my_rom(12699);
when "00111111001" => 
 data1 <= my_rom(505); 
 data2 <= my_rom(1860); 
 data3 <= my_rom(3215); 
 data4 <= my_rom(4570); 
 data5 <= my_rom(5925); 
 data6 <= my_rom(7280); 
 data7 <= my_rom(8635); 
 data8 <= my_rom(9990); 
 data9 <= my_rom(11345); 
 data10 <= my_rom(12700);
when "00111111010" => 
 data1 <= my_rom(506); 
 data2 <= my_rom(1861); 
 data3 <= my_rom(3216); 
 data4 <= my_rom(4571); 
 data5 <= my_rom(5926); 
 data6 <= my_rom(7281); 
 data7 <= my_rom(8636); 
 data8 <= my_rom(9991); 
 data9 <= my_rom(11346); 
 data10 <= my_rom(12701);
when "00111111011" => 
 data1 <= my_rom(507); 
 data2 <= my_rom(1862); 
 data3 <= my_rom(3217); 
 data4 <= my_rom(4572); 
 data5 <= my_rom(5927); 
 data6 <= my_rom(7282); 
 data7 <= my_rom(8637); 
 data8 <= my_rom(9992); 
 data9 <= my_rom(11347); 
 data10 <= my_rom(12702);
when "00111111100" => 
 data1 <= my_rom(508); 
 data2 <= my_rom(1863); 
 data3 <= my_rom(3218); 
 data4 <= my_rom(4573); 
 data5 <= my_rom(5928); 
 data6 <= my_rom(7283); 
 data7 <= my_rom(8638); 
 data8 <= my_rom(9993); 
 data9 <= my_rom(11348); 
 data10 <= my_rom(12703);
when "00111111101" => 
 data1 <= my_rom(509); 
 data2 <= my_rom(1864); 
 data3 <= my_rom(3219); 
 data4 <= my_rom(4574); 
 data5 <= my_rom(5929); 
 data6 <= my_rom(7284); 
 data7 <= my_rom(8639); 
 data8 <= my_rom(9994); 
 data9 <= my_rom(11349); 
 data10 <= my_rom(12704);
when "00111111110" => 
 data1 <= my_rom(510); 
 data2 <= my_rom(1865); 
 data3 <= my_rom(3220); 
 data4 <= my_rom(4575); 
 data5 <= my_rom(5930); 
 data6 <= my_rom(7285); 
 data7 <= my_rom(8640); 
 data8 <= my_rom(9995); 
 data9 <= my_rom(11350); 
 data10 <= my_rom(12705);
when "00111111111" => 
 data1 <= my_rom(511); 
 data2 <= my_rom(1866); 
 data3 <= my_rom(3221); 
 data4 <= my_rom(4576); 
 data5 <= my_rom(5931); 
 data6 <= my_rom(7286); 
 data7 <= my_rom(8641); 
 data8 <= my_rom(9996); 
 data9 <= my_rom(11351); 
 data10 <= my_rom(12706);
when "01000000000" => 
 data1 <= my_rom(512); 
 data2 <= my_rom(1867); 
 data3 <= my_rom(3222); 
 data4 <= my_rom(4577); 
 data5 <= my_rom(5932); 
 data6 <= my_rom(7287); 
 data7 <= my_rom(8642); 
 data8 <= my_rom(9997); 
 data9 <= my_rom(11352); 
 data10 <= my_rom(12707);
when "01000000001" => 
 data1 <= my_rom(513); 
 data2 <= my_rom(1868); 
 data3 <= my_rom(3223); 
 data4 <= my_rom(4578); 
 data5 <= my_rom(5933); 
 data6 <= my_rom(7288); 
 data7 <= my_rom(8643); 
 data8 <= my_rom(9998); 
 data9 <= my_rom(11353); 
 data10 <= my_rom(12708);
when "01000000010" => 
 data1 <= my_rom(514); 
 data2 <= my_rom(1869); 
 data3 <= my_rom(3224); 
 data4 <= my_rom(4579); 
 data5 <= my_rom(5934); 
 data6 <= my_rom(7289); 
 data7 <= my_rom(8644); 
 data8 <= my_rom(9999); 
 data9 <= my_rom(11354); 
 data10 <= my_rom(12709);
when "01000000011" => 
 data1 <= my_rom(515); 
 data2 <= my_rom(1870); 
 data3 <= my_rom(3225); 
 data4 <= my_rom(4580); 
 data5 <= my_rom(5935); 
 data6 <= my_rom(7290); 
 data7 <= my_rom(8645); 
 data8 <= my_rom(10000); 
 data9 <= my_rom(11355); 
 data10 <= my_rom(12710);
when "01000000100" => 
 data1 <= my_rom(516); 
 data2 <= my_rom(1871); 
 data3 <= my_rom(3226); 
 data4 <= my_rom(4581); 
 data5 <= my_rom(5936); 
 data6 <= my_rom(7291); 
 data7 <= my_rom(8646); 
 data8 <= my_rom(10001); 
 data9 <= my_rom(11356); 
 data10 <= my_rom(12711);
when "01000000101" => 
 data1 <= my_rom(517); 
 data2 <= my_rom(1872); 
 data3 <= my_rom(3227); 
 data4 <= my_rom(4582); 
 data5 <= my_rom(5937); 
 data6 <= my_rom(7292); 
 data7 <= my_rom(8647); 
 data8 <= my_rom(10002); 
 data9 <= my_rom(11357); 
 data10 <= my_rom(12712);
when "01000000110" => 
 data1 <= my_rom(518); 
 data2 <= my_rom(1873); 
 data3 <= my_rom(3228); 
 data4 <= my_rom(4583); 
 data5 <= my_rom(5938); 
 data6 <= my_rom(7293); 
 data7 <= my_rom(8648); 
 data8 <= my_rom(10003); 
 data9 <= my_rom(11358); 
 data10 <= my_rom(12713);
when "01000000111" => 
 data1 <= my_rom(519); 
 data2 <= my_rom(1874); 
 data3 <= my_rom(3229); 
 data4 <= my_rom(4584); 
 data5 <= my_rom(5939); 
 data6 <= my_rom(7294); 
 data7 <= my_rom(8649); 
 data8 <= my_rom(10004); 
 data9 <= my_rom(11359); 
 data10 <= my_rom(12714);
when "01000001000" => 
 data1 <= my_rom(520); 
 data2 <= my_rom(1875); 
 data3 <= my_rom(3230); 
 data4 <= my_rom(4585); 
 data5 <= my_rom(5940); 
 data6 <= my_rom(7295); 
 data7 <= my_rom(8650); 
 data8 <= my_rom(10005); 
 data9 <= my_rom(11360); 
 data10 <= my_rom(12715);
when "01000001001" => 
 data1 <= my_rom(521); 
 data2 <= my_rom(1876); 
 data3 <= my_rom(3231); 
 data4 <= my_rom(4586); 
 data5 <= my_rom(5941); 
 data6 <= my_rom(7296); 
 data7 <= my_rom(8651); 
 data8 <= my_rom(10006); 
 data9 <= my_rom(11361); 
 data10 <= my_rom(12716);
when "01000001010" => 
 data1 <= my_rom(522); 
 data2 <= my_rom(1877); 
 data3 <= my_rom(3232); 
 data4 <= my_rom(4587); 
 data5 <= my_rom(5942); 
 data6 <= my_rom(7297); 
 data7 <= my_rom(8652); 
 data8 <= my_rom(10007); 
 data9 <= my_rom(11362); 
 data10 <= my_rom(12717);
when "01000001011" => 
 data1 <= my_rom(523); 
 data2 <= my_rom(1878); 
 data3 <= my_rom(3233); 
 data4 <= my_rom(4588); 
 data5 <= my_rom(5943); 
 data6 <= my_rom(7298); 
 data7 <= my_rom(8653); 
 data8 <= my_rom(10008); 
 data9 <= my_rom(11363); 
 data10 <= my_rom(12718);
when "01000001100" => 
 data1 <= my_rom(524); 
 data2 <= my_rom(1879); 
 data3 <= my_rom(3234); 
 data4 <= my_rom(4589); 
 data5 <= my_rom(5944); 
 data6 <= my_rom(7299); 
 data7 <= my_rom(8654); 
 data8 <= my_rom(10009); 
 data9 <= my_rom(11364); 
 data10 <= my_rom(12719);
when "01000001101" => 
 data1 <= my_rom(525); 
 data2 <= my_rom(1880); 
 data3 <= my_rom(3235); 
 data4 <= my_rom(4590); 
 data5 <= my_rom(5945); 
 data6 <= my_rom(7300); 
 data7 <= my_rom(8655); 
 data8 <= my_rom(10010); 
 data9 <= my_rom(11365); 
 data10 <= my_rom(12720);
when "01000001110" => 
 data1 <= my_rom(526); 
 data2 <= my_rom(1881); 
 data3 <= my_rom(3236); 
 data4 <= my_rom(4591); 
 data5 <= my_rom(5946); 
 data6 <= my_rom(7301); 
 data7 <= my_rom(8656); 
 data8 <= my_rom(10011); 
 data9 <= my_rom(11366); 
 data10 <= my_rom(12721);
when "01000001111" => 
 data1 <= my_rom(527); 
 data2 <= my_rom(1882); 
 data3 <= my_rom(3237); 
 data4 <= my_rom(4592); 
 data5 <= my_rom(5947); 
 data6 <= my_rom(7302); 
 data7 <= my_rom(8657); 
 data8 <= my_rom(10012); 
 data9 <= my_rom(11367); 
 data10 <= my_rom(12722);
when "01000010000" => 
 data1 <= my_rom(528); 
 data2 <= my_rom(1883); 
 data3 <= my_rom(3238); 
 data4 <= my_rom(4593); 
 data5 <= my_rom(5948); 
 data6 <= my_rom(7303); 
 data7 <= my_rom(8658); 
 data8 <= my_rom(10013); 
 data9 <= my_rom(11368); 
 data10 <= my_rom(12723);
when "01000010001" => 
 data1 <= my_rom(529); 
 data2 <= my_rom(1884); 
 data3 <= my_rom(3239); 
 data4 <= my_rom(4594); 
 data5 <= my_rom(5949); 
 data6 <= my_rom(7304); 
 data7 <= my_rom(8659); 
 data8 <= my_rom(10014); 
 data9 <= my_rom(11369); 
 data10 <= my_rom(12724);
when "01000010010" => 
 data1 <= my_rom(530); 
 data2 <= my_rom(1885); 
 data3 <= my_rom(3240); 
 data4 <= my_rom(4595); 
 data5 <= my_rom(5950); 
 data6 <= my_rom(7305); 
 data7 <= my_rom(8660); 
 data8 <= my_rom(10015); 
 data9 <= my_rom(11370); 
 data10 <= my_rom(12725);
when "01000010011" => 
 data1 <= my_rom(531); 
 data2 <= my_rom(1886); 
 data3 <= my_rom(3241); 
 data4 <= my_rom(4596); 
 data5 <= my_rom(5951); 
 data6 <= my_rom(7306); 
 data7 <= my_rom(8661); 
 data8 <= my_rom(10016); 
 data9 <= my_rom(11371); 
 data10 <= my_rom(12726);
when "01000010100" => 
 data1 <= my_rom(532); 
 data2 <= my_rom(1887); 
 data3 <= my_rom(3242); 
 data4 <= my_rom(4597); 
 data5 <= my_rom(5952); 
 data6 <= my_rom(7307); 
 data7 <= my_rom(8662); 
 data8 <= my_rom(10017); 
 data9 <= my_rom(11372); 
 data10 <= my_rom(12727);
when "01000010101" => 
 data1 <= my_rom(533); 
 data2 <= my_rom(1888); 
 data3 <= my_rom(3243); 
 data4 <= my_rom(4598); 
 data5 <= my_rom(5953); 
 data6 <= my_rom(7308); 
 data7 <= my_rom(8663); 
 data8 <= my_rom(10018); 
 data9 <= my_rom(11373); 
 data10 <= my_rom(12728);
when "01000010110" => 
 data1 <= my_rom(534); 
 data2 <= my_rom(1889); 
 data3 <= my_rom(3244); 
 data4 <= my_rom(4599); 
 data5 <= my_rom(5954); 
 data6 <= my_rom(7309); 
 data7 <= my_rom(8664); 
 data8 <= my_rom(10019); 
 data9 <= my_rom(11374); 
 data10 <= my_rom(12729);
when "01000010111" => 
 data1 <= my_rom(535); 
 data2 <= my_rom(1890); 
 data3 <= my_rom(3245); 
 data4 <= my_rom(4600); 
 data5 <= my_rom(5955); 
 data6 <= my_rom(7310); 
 data7 <= my_rom(8665); 
 data8 <= my_rom(10020); 
 data9 <= my_rom(11375); 
 data10 <= my_rom(12730);
when "01000011000" => 
 data1 <= my_rom(536); 
 data2 <= my_rom(1891); 
 data3 <= my_rom(3246); 
 data4 <= my_rom(4601); 
 data5 <= my_rom(5956); 
 data6 <= my_rom(7311); 
 data7 <= my_rom(8666); 
 data8 <= my_rom(10021); 
 data9 <= my_rom(11376); 
 data10 <= my_rom(12731);
when "01000011001" => 
 data1 <= my_rom(537); 
 data2 <= my_rom(1892); 
 data3 <= my_rom(3247); 
 data4 <= my_rom(4602); 
 data5 <= my_rom(5957); 
 data6 <= my_rom(7312); 
 data7 <= my_rom(8667); 
 data8 <= my_rom(10022); 
 data9 <= my_rom(11377); 
 data10 <= my_rom(12732);
when "01000011010" => 
 data1 <= my_rom(538); 
 data2 <= my_rom(1893); 
 data3 <= my_rom(3248); 
 data4 <= my_rom(4603); 
 data5 <= my_rom(5958); 
 data6 <= my_rom(7313); 
 data7 <= my_rom(8668); 
 data8 <= my_rom(10023); 
 data9 <= my_rom(11378); 
 data10 <= my_rom(12733);
when "01000011011" => 
 data1 <= my_rom(539); 
 data2 <= my_rom(1894); 
 data3 <= my_rom(3249); 
 data4 <= my_rom(4604); 
 data5 <= my_rom(5959); 
 data6 <= my_rom(7314); 
 data7 <= my_rom(8669); 
 data8 <= my_rom(10024); 
 data9 <= my_rom(11379); 
 data10 <= my_rom(12734);
when "01000011100" => 
 data1 <= my_rom(540); 
 data2 <= my_rom(1895); 
 data3 <= my_rom(3250); 
 data4 <= my_rom(4605); 
 data5 <= my_rom(5960); 
 data6 <= my_rom(7315); 
 data7 <= my_rom(8670); 
 data8 <= my_rom(10025); 
 data9 <= my_rom(11380); 
 data10 <= my_rom(12735);
when "01000011101" => 
 data1 <= my_rom(541); 
 data2 <= my_rom(1896); 
 data3 <= my_rom(3251); 
 data4 <= my_rom(4606); 
 data5 <= my_rom(5961); 
 data6 <= my_rom(7316); 
 data7 <= my_rom(8671); 
 data8 <= my_rom(10026); 
 data9 <= my_rom(11381); 
 data10 <= my_rom(12736);
when "01000011110" => 
 data1 <= my_rom(542); 
 data2 <= my_rom(1897); 
 data3 <= my_rom(3252); 
 data4 <= my_rom(4607); 
 data5 <= my_rom(5962); 
 data6 <= my_rom(7317); 
 data7 <= my_rom(8672); 
 data8 <= my_rom(10027); 
 data9 <= my_rom(11382); 
 data10 <= my_rom(12737);
when "01000011111" => 
 data1 <= my_rom(543); 
 data2 <= my_rom(1898); 
 data3 <= my_rom(3253); 
 data4 <= my_rom(4608); 
 data5 <= my_rom(5963); 
 data6 <= my_rom(7318); 
 data7 <= my_rom(8673); 
 data8 <= my_rom(10028); 
 data9 <= my_rom(11383); 
 data10 <= my_rom(12738);
when "01000100000" => 
 data1 <= my_rom(544); 
 data2 <= my_rom(1899); 
 data3 <= my_rom(3254); 
 data4 <= my_rom(4609); 
 data5 <= my_rom(5964); 
 data6 <= my_rom(7319); 
 data7 <= my_rom(8674); 
 data8 <= my_rom(10029); 
 data9 <= my_rom(11384); 
 data10 <= my_rom(12739);
when "01000100001" => 
 data1 <= my_rom(545); 
 data2 <= my_rom(1900); 
 data3 <= my_rom(3255); 
 data4 <= my_rom(4610); 
 data5 <= my_rom(5965); 
 data6 <= my_rom(7320); 
 data7 <= my_rom(8675); 
 data8 <= my_rom(10030); 
 data9 <= my_rom(11385); 
 data10 <= my_rom(12740);
when "01000100010" => 
 data1 <= my_rom(546); 
 data2 <= my_rom(1901); 
 data3 <= my_rom(3256); 
 data4 <= my_rom(4611); 
 data5 <= my_rom(5966); 
 data6 <= my_rom(7321); 
 data7 <= my_rom(8676); 
 data8 <= my_rom(10031); 
 data9 <= my_rom(11386); 
 data10 <= my_rom(12741);
when "01000100011" => 
 data1 <= my_rom(547); 
 data2 <= my_rom(1902); 
 data3 <= my_rom(3257); 
 data4 <= my_rom(4612); 
 data5 <= my_rom(5967); 
 data6 <= my_rom(7322); 
 data7 <= my_rom(8677); 
 data8 <= my_rom(10032); 
 data9 <= my_rom(11387); 
 data10 <= my_rom(12742);
when "01000100100" => 
 data1 <= my_rom(548); 
 data2 <= my_rom(1903); 
 data3 <= my_rom(3258); 
 data4 <= my_rom(4613); 
 data5 <= my_rom(5968); 
 data6 <= my_rom(7323); 
 data7 <= my_rom(8678); 
 data8 <= my_rom(10033); 
 data9 <= my_rom(11388); 
 data10 <= my_rom(12743);
when "01000100101" => 
 data1 <= my_rom(549); 
 data2 <= my_rom(1904); 
 data3 <= my_rom(3259); 
 data4 <= my_rom(4614); 
 data5 <= my_rom(5969); 
 data6 <= my_rom(7324); 
 data7 <= my_rom(8679); 
 data8 <= my_rom(10034); 
 data9 <= my_rom(11389); 
 data10 <= my_rom(12744);
when "01000100110" => 
 data1 <= my_rom(550); 
 data2 <= my_rom(1905); 
 data3 <= my_rom(3260); 
 data4 <= my_rom(4615); 
 data5 <= my_rom(5970); 
 data6 <= my_rom(7325); 
 data7 <= my_rom(8680); 
 data8 <= my_rom(10035); 
 data9 <= my_rom(11390); 
 data10 <= my_rom(12745);
when "01000100111" => 
 data1 <= my_rom(551); 
 data2 <= my_rom(1906); 
 data3 <= my_rom(3261); 
 data4 <= my_rom(4616); 
 data5 <= my_rom(5971); 
 data6 <= my_rom(7326); 
 data7 <= my_rom(8681); 
 data8 <= my_rom(10036); 
 data9 <= my_rom(11391); 
 data10 <= my_rom(12746);
when "01000101000" => 
 data1 <= my_rom(552); 
 data2 <= my_rom(1907); 
 data3 <= my_rom(3262); 
 data4 <= my_rom(4617); 
 data5 <= my_rom(5972); 
 data6 <= my_rom(7327); 
 data7 <= my_rom(8682); 
 data8 <= my_rom(10037); 
 data9 <= my_rom(11392); 
 data10 <= my_rom(12747);
when "01000101001" => 
 data1 <= my_rom(553); 
 data2 <= my_rom(1908); 
 data3 <= my_rom(3263); 
 data4 <= my_rom(4618); 
 data5 <= my_rom(5973); 
 data6 <= my_rom(7328); 
 data7 <= my_rom(8683); 
 data8 <= my_rom(10038); 
 data9 <= my_rom(11393); 
 data10 <= my_rom(12748);
when "01000101010" => 
 data1 <= my_rom(554); 
 data2 <= my_rom(1909); 
 data3 <= my_rom(3264); 
 data4 <= my_rom(4619); 
 data5 <= my_rom(5974); 
 data6 <= my_rom(7329); 
 data7 <= my_rom(8684); 
 data8 <= my_rom(10039); 
 data9 <= my_rom(11394); 
 data10 <= my_rom(12749);
when "01000101011" => 
 data1 <= my_rom(555); 
 data2 <= my_rom(1910); 
 data3 <= my_rom(3265); 
 data4 <= my_rom(4620); 
 data5 <= my_rom(5975); 
 data6 <= my_rom(7330); 
 data7 <= my_rom(8685); 
 data8 <= my_rom(10040); 
 data9 <= my_rom(11395); 
 data10 <= my_rom(12750);
when "01000101100" => 
 data1 <= my_rom(556); 
 data2 <= my_rom(1911); 
 data3 <= my_rom(3266); 
 data4 <= my_rom(4621); 
 data5 <= my_rom(5976); 
 data6 <= my_rom(7331); 
 data7 <= my_rom(8686); 
 data8 <= my_rom(10041); 
 data9 <= my_rom(11396); 
 data10 <= my_rom(12751);
when "01000101101" => 
 data1 <= my_rom(557); 
 data2 <= my_rom(1912); 
 data3 <= my_rom(3267); 
 data4 <= my_rom(4622); 
 data5 <= my_rom(5977); 
 data6 <= my_rom(7332); 
 data7 <= my_rom(8687); 
 data8 <= my_rom(10042); 
 data9 <= my_rom(11397); 
 data10 <= my_rom(12752);
when "01000101110" => 
 data1 <= my_rom(558); 
 data2 <= my_rom(1913); 
 data3 <= my_rom(3268); 
 data4 <= my_rom(4623); 
 data5 <= my_rom(5978); 
 data6 <= my_rom(7333); 
 data7 <= my_rom(8688); 
 data8 <= my_rom(10043); 
 data9 <= my_rom(11398); 
 data10 <= my_rom(12753);
when "01000101111" => 
 data1 <= my_rom(559); 
 data2 <= my_rom(1914); 
 data3 <= my_rom(3269); 
 data4 <= my_rom(4624); 
 data5 <= my_rom(5979); 
 data6 <= my_rom(7334); 
 data7 <= my_rom(8689); 
 data8 <= my_rom(10044); 
 data9 <= my_rom(11399); 
 data10 <= my_rom(12754);
when "01000110000" => 
 data1 <= my_rom(560); 
 data2 <= my_rom(1915); 
 data3 <= my_rom(3270); 
 data4 <= my_rom(4625); 
 data5 <= my_rom(5980); 
 data6 <= my_rom(7335); 
 data7 <= my_rom(8690); 
 data8 <= my_rom(10045); 
 data9 <= my_rom(11400); 
 data10 <= my_rom(12755);
when "01000110001" => 
 data1 <= my_rom(561); 
 data2 <= my_rom(1916); 
 data3 <= my_rom(3271); 
 data4 <= my_rom(4626); 
 data5 <= my_rom(5981); 
 data6 <= my_rom(7336); 
 data7 <= my_rom(8691); 
 data8 <= my_rom(10046); 
 data9 <= my_rom(11401); 
 data10 <= my_rom(12756);
when "01000110010" => 
 data1 <= my_rom(562); 
 data2 <= my_rom(1917); 
 data3 <= my_rom(3272); 
 data4 <= my_rom(4627); 
 data5 <= my_rom(5982); 
 data6 <= my_rom(7337); 
 data7 <= my_rom(8692); 
 data8 <= my_rom(10047); 
 data9 <= my_rom(11402); 
 data10 <= my_rom(12757);
when "01000110011" => 
 data1 <= my_rom(563); 
 data2 <= my_rom(1918); 
 data3 <= my_rom(3273); 
 data4 <= my_rom(4628); 
 data5 <= my_rom(5983); 
 data6 <= my_rom(7338); 
 data7 <= my_rom(8693); 
 data8 <= my_rom(10048); 
 data9 <= my_rom(11403); 
 data10 <= my_rom(12758);
when "01000110100" => 
 data1 <= my_rom(564); 
 data2 <= my_rom(1919); 
 data3 <= my_rom(3274); 
 data4 <= my_rom(4629); 
 data5 <= my_rom(5984); 
 data6 <= my_rom(7339); 
 data7 <= my_rom(8694); 
 data8 <= my_rom(10049); 
 data9 <= my_rom(11404); 
 data10 <= my_rom(12759);
when "01000110101" => 
 data1 <= my_rom(565); 
 data2 <= my_rom(1920); 
 data3 <= my_rom(3275); 
 data4 <= my_rom(4630); 
 data5 <= my_rom(5985); 
 data6 <= my_rom(7340); 
 data7 <= my_rom(8695); 
 data8 <= my_rom(10050); 
 data9 <= my_rom(11405); 
 data10 <= my_rom(12760);
when "01000110110" => 
 data1 <= my_rom(566); 
 data2 <= my_rom(1921); 
 data3 <= my_rom(3276); 
 data4 <= my_rom(4631); 
 data5 <= my_rom(5986); 
 data6 <= my_rom(7341); 
 data7 <= my_rom(8696); 
 data8 <= my_rom(10051); 
 data9 <= my_rom(11406); 
 data10 <= my_rom(12761);
when "01000110111" => 
 data1 <= my_rom(567); 
 data2 <= my_rom(1922); 
 data3 <= my_rom(3277); 
 data4 <= my_rom(4632); 
 data5 <= my_rom(5987); 
 data6 <= my_rom(7342); 
 data7 <= my_rom(8697); 
 data8 <= my_rom(10052); 
 data9 <= my_rom(11407); 
 data10 <= my_rom(12762);
when "01000111000" => 
 data1 <= my_rom(568); 
 data2 <= my_rom(1923); 
 data3 <= my_rom(3278); 
 data4 <= my_rom(4633); 
 data5 <= my_rom(5988); 
 data6 <= my_rom(7343); 
 data7 <= my_rom(8698); 
 data8 <= my_rom(10053); 
 data9 <= my_rom(11408); 
 data10 <= my_rom(12763);
when "01000111001" => 
 data1 <= my_rom(569); 
 data2 <= my_rom(1924); 
 data3 <= my_rom(3279); 
 data4 <= my_rom(4634); 
 data5 <= my_rom(5989); 
 data6 <= my_rom(7344); 
 data7 <= my_rom(8699); 
 data8 <= my_rom(10054); 
 data9 <= my_rom(11409); 
 data10 <= my_rom(12764);
when "01000111010" => 
 data1 <= my_rom(570); 
 data2 <= my_rom(1925); 
 data3 <= my_rom(3280); 
 data4 <= my_rom(4635); 
 data5 <= my_rom(5990); 
 data6 <= my_rom(7345); 
 data7 <= my_rom(8700); 
 data8 <= my_rom(10055); 
 data9 <= my_rom(11410); 
 data10 <= my_rom(12765);
when "01000111011" => 
 data1 <= my_rom(571); 
 data2 <= my_rom(1926); 
 data3 <= my_rom(3281); 
 data4 <= my_rom(4636); 
 data5 <= my_rom(5991); 
 data6 <= my_rom(7346); 
 data7 <= my_rom(8701); 
 data8 <= my_rom(10056); 
 data9 <= my_rom(11411); 
 data10 <= my_rom(12766);
when "01000111100" => 
 data1 <= my_rom(572); 
 data2 <= my_rom(1927); 
 data3 <= my_rom(3282); 
 data4 <= my_rom(4637); 
 data5 <= my_rom(5992); 
 data6 <= my_rom(7347); 
 data7 <= my_rom(8702); 
 data8 <= my_rom(10057); 
 data9 <= my_rom(11412); 
 data10 <= my_rom(12767);
when "01000111101" => 
 data1 <= my_rom(573); 
 data2 <= my_rom(1928); 
 data3 <= my_rom(3283); 
 data4 <= my_rom(4638); 
 data5 <= my_rom(5993); 
 data6 <= my_rom(7348); 
 data7 <= my_rom(8703); 
 data8 <= my_rom(10058); 
 data9 <= my_rom(11413); 
 data10 <= my_rom(12768);
when "01000111110" => 
 data1 <= my_rom(574); 
 data2 <= my_rom(1929); 
 data3 <= my_rom(3284); 
 data4 <= my_rom(4639); 
 data5 <= my_rom(5994); 
 data6 <= my_rom(7349); 
 data7 <= my_rom(8704); 
 data8 <= my_rom(10059); 
 data9 <= my_rom(11414); 
 data10 <= my_rom(12769);
when "01000111111" => 
 data1 <= my_rom(575); 
 data2 <= my_rom(1930); 
 data3 <= my_rom(3285); 
 data4 <= my_rom(4640); 
 data5 <= my_rom(5995); 
 data6 <= my_rom(7350); 
 data7 <= my_rom(8705); 
 data8 <= my_rom(10060); 
 data9 <= my_rom(11415); 
 data10 <= my_rom(12770);
when "01001000000" => 
 data1 <= my_rom(576); 
 data2 <= my_rom(1931); 
 data3 <= my_rom(3286); 
 data4 <= my_rom(4641); 
 data5 <= my_rom(5996); 
 data6 <= my_rom(7351); 
 data7 <= my_rom(8706); 
 data8 <= my_rom(10061); 
 data9 <= my_rom(11416); 
 data10 <= my_rom(12771);
when "01001000001" => 
 data1 <= my_rom(577); 
 data2 <= my_rom(1932); 
 data3 <= my_rom(3287); 
 data4 <= my_rom(4642); 
 data5 <= my_rom(5997); 
 data6 <= my_rom(7352); 
 data7 <= my_rom(8707); 
 data8 <= my_rom(10062); 
 data9 <= my_rom(11417); 
 data10 <= my_rom(12772);
when "01001000010" => 
 data1 <= my_rom(578); 
 data2 <= my_rom(1933); 
 data3 <= my_rom(3288); 
 data4 <= my_rom(4643); 
 data5 <= my_rom(5998); 
 data6 <= my_rom(7353); 
 data7 <= my_rom(8708); 
 data8 <= my_rom(10063); 
 data9 <= my_rom(11418); 
 data10 <= my_rom(12773);
when "01001000011" => 
 data1 <= my_rom(579); 
 data2 <= my_rom(1934); 
 data3 <= my_rom(3289); 
 data4 <= my_rom(4644); 
 data5 <= my_rom(5999); 
 data6 <= my_rom(7354); 
 data7 <= my_rom(8709); 
 data8 <= my_rom(10064); 
 data9 <= my_rom(11419); 
 data10 <= my_rom(12774);
when "01001000100" => 
 data1 <= my_rom(580); 
 data2 <= my_rom(1935); 
 data3 <= my_rom(3290); 
 data4 <= my_rom(4645); 
 data5 <= my_rom(6000); 
 data6 <= my_rom(7355); 
 data7 <= my_rom(8710); 
 data8 <= my_rom(10065); 
 data9 <= my_rom(11420); 
 data10 <= my_rom(12775);
when "01001000101" => 
 data1 <= my_rom(581); 
 data2 <= my_rom(1936); 
 data3 <= my_rom(3291); 
 data4 <= my_rom(4646); 
 data5 <= my_rom(6001); 
 data6 <= my_rom(7356); 
 data7 <= my_rom(8711); 
 data8 <= my_rom(10066); 
 data9 <= my_rom(11421); 
 data10 <= my_rom(12776);
when "01001000110" => 
 data1 <= my_rom(582); 
 data2 <= my_rom(1937); 
 data3 <= my_rom(3292); 
 data4 <= my_rom(4647); 
 data5 <= my_rom(6002); 
 data6 <= my_rom(7357); 
 data7 <= my_rom(8712); 
 data8 <= my_rom(10067); 
 data9 <= my_rom(11422); 
 data10 <= my_rom(12777);
when "01001000111" => 
 data1 <= my_rom(583); 
 data2 <= my_rom(1938); 
 data3 <= my_rom(3293); 
 data4 <= my_rom(4648); 
 data5 <= my_rom(6003); 
 data6 <= my_rom(7358); 
 data7 <= my_rom(8713); 
 data8 <= my_rom(10068); 
 data9 <= my_rom(11423); 
 data10 <= my_rom(12778);
when "01001001000" => 
 data1 <= my_rom(584); 
 data2 <= my_rom(1939); 
 data3 <= my_rom(3294); 
 data4 <= my_rom(4649); 
 data5 <= my_rom(6004); 
 data6 <= my_rom(7359); 
 data7 <= my_rom(8714); 
 data8 <= my_rom(10069); 
 data9 <= my_rom(11424); 
 data10 <= my_rom(12779);
when "01001001001" => 
 data1 <= my_rom(585); 
 data2 <= my_rom(1940); 
 data3 <= my_rom(3295); 
 data4 <= my_rom(4650); 
 data5 <= my_rom(6005); 
 data6 <= my_rom(7360); 
 data7 <= my_rom(8715); 
 data8 <= my_rom(10070); 
 data9 <= my_rom(11425); 
 data10 <= my_rom(12780);
when "01001001010" => 
 data1 <= my_rom(586); 
 data2 <= my_rom(1941); 
 data3 <= my_rom(3296); 
 data4 <= my_rom(4651); 
 data5 <= my_rom(6006); 
 data6 <= my_rom(7361); 
 data7 <= my_rom(8716); 
 data8 <= my_rom(10071); 
 data9 <= my_rom(11426); 
 data10 <= my_rom(12781);
when "01001001011" => 
 data1 <= my_rom(587); 
 data2 <= my_rom(1942); 
 data3 <= my_rom(3297); 
 data4 <= my_rom(4652); 
 data5 <= my_rom(6007); 
 data6 <= my_rom(7362); 
 data7 <= my_rom(8717); 
 data8 <= my_rom(10072); 
 data9 <= my_rom(11427); 
 data10 <= my_rom(12782);
when "01001001100" => 
 data1 <= my_rom(588); 
 data2 <= my_rom(1943); 
 data3 <= my_rom(3298); 
 data4 <= my_rom(4653); 
 data5 <= my_rom(6008); 
 data6 <= my_rom(7363); 
 data7 <= my_rom(8718); 
 data8 <= my_rom(10073); 
 data9 <= my_rom(11428); 
 data10 <= my_rom(12783);
when "01001001101" => 
 data1 <= my_rom(589); 
 data2 <= my_rom(1944); 
 data3 <= my_rom(3299); 
 data4 <= my_rom(4654); 
 data5 <= my_rom(6009); 
 data6 <= my_rom(7364); 
 data7 <= my_rom(8719); 
 data8 <= my_rom(10074); 
 data9 <= my_rom(11429); 
 data10 <= my_rom(12784);
when "01001001110" => 
 data1 <= my_rom(590); 
 data2 <= my_rom(1945); 
 data3 <= my_rom(3300); 
 data4 <= my_rom(4655); 
 data5 <= my_rom(6010); 
 data6 <= my_rom(7365); 
 data7 <= my_rom(8720); 
 data8 <= my_rom(10075); 
 data9 <= my_rom(11430); 
 data10 <= my_rom(12785);
when "01001001111" => 
 data1 <= my_rom(591); 
 data2 <= my_rom(1946); 
 data3 <= my_rom(3301); 
 data4 <= my_rom(4656); 
 data5 <= my_rom(6011); 
 data6 <= my_rom(7366); 
 data7 <= my_rom(8721); 
 data8 <= my_rom(10076); 
 data9 <= my_rom(11431); 
 data10 <= my_rom(12786);
when "01001010000" => 
 data1 <= my_rom(592); 
 data2 <= my_rom(1947); 
 data3 <= my_rom(3302); 
 data4 <= my_rom(4657); 
 data5 <= my_rom(6012); 
 data6 <= my_rom(7367); 
 data7 <= my_rom(8722); 
 data8 <= my_rom(10077); 
 data9 <= my_rom(11432); 
 data10 <= my_rom(12787);
when "01001010001" => 
 data1 <= my_rom(593); 
 data2 <= my_rom(1948); 
 data3 <= my_rom(3303); 
 data4 <= my_rom(4658); 
 data5 <= my_rom(6013); 
 data6 <= my_rom(7368); 
 data7 <= my_rom(8723); 
 data8 <= my_rom(10078); 
 data9 <= my_rom(11433); 
 data10 <= my_rom(12788);
when "01001010010" => 
 data1 <= my_rom(594); 
 data2 <= my_rom(1949); 
 data3 <= my_rom(3304); 
 data4 <= my_rom(4659); 
 data5 <= my_rom(6014); 
 data6 <= my_rom(7369); 
 data7 <= my_rom(8724); 
 data8 <= my_rom(10079); 
 data9 <= my_rom(11434); 
 data10 <= my_rom(12789);
when "01001010011" => 
 data1 <= my_rom(595); 
 data2 <= my_rom(1950); 
 data3 <= my_rom(3305); 
 data4 <= my_rom(4660); 
 data5 <= my_rom(6015); 
 data6 <= my_rom(7370); 
 data7 <= my_rom(8725); 
 data8 <= my_rom(10080); 
 data9 <= my_rom(11435); 
 data10 <= my_rom(12790);
when "01001010100" => 
 data1 <= my_rom(596); 
 data2 <= my_rom(1951); 
 data3 <= my_rom(3306); 
 data4 <= my_rom(4661); 
 data5 <= my_rom(6016); 
 data6 <= my_rom(7371); 
 data7 <= my_rom(8726); 
 data8 <= my_rom(10081); 
 data9 <= my_rom(11436); 
 data10 <= my_rom(12791);
when "01001010101" => 
 data1 <= my_rom(597); 
 data2 <= my_rom(1952); 
 data3 <= my_rom(3307); 
 data4 <= my_rom(4662); 
 data5 <= my_rom(6017); 
 data6 <= my_rom(7372); 
 data7 <= my_rom(8727); 
 data8 <= my_rom(10082); 
 data9 <= my_rom(11437); 
 data10 <= my_rom(12792);
when "01001010110" => 
 data1 <= my_rom(598); 
 data2 <= my_rom(1953); 
 data3 <= my_rom(3308); 
 data4 <= my_rom(4663); 
 data5 <= my_rom(6018); 
 data6 <= my_rom(7373); 
 data7 <= my_rom(8728); 
 data8 <= my_rom(10083); 
 data9 <= my_rom(11438); 
 data10 <= my_rom(12793);
when "01001010111" => 
 data1 <= my_rom(599); 
 data2 <= my_rom(1954); 
 data3 <= my_rom(3309); 
 data4 <= my_rom(4664); 
 data5 <= my_rom(6019); 
 data6 <= my_rom(7374); 
 data7 <= my_rom(8729); 
 data8 <= my_rom(10084); 
 data9 <= my_rom(11439); 
 data10 <= my_rom(12794);
when "01001011000" => 
 data1 <= my_rom(600); 
 data2 <= my_rom(1955); 
 data3 <= my_rom(3310); 
 data4 <= my_rom(4665); 
 data5 <= my_rom(6020); 
 data6 <= my_rom(7375); 
 data7 <= my_rom(8730); 
 data8 <= my_rom(10085); 
 data9 <= my_rom(11440); 
 data10 <= my_rom(12795);
when "01001011001" => 
 data1 <= my_rom(601); 
 data2 <= my_rom(1956); 
 data3 <= my_rom(3311); 
 data4 <= my_rom(4666); 
 data5 <= my_rom(6021); 
 data6 <= my_rom(7376); 
 data7 <= my_rom(8731); 
 data8 <= my_rom(10086); 
 data9 <= my_rom(11441); 
 data10 <= my_rom(12796);
when "01001011010" => 
 data1 <= my_rom(602); 
 data2 <= my_rom(1957); 
 data3 <= my_rom(3312); 
 data4 <= my_rom(4667); 
 data5 <= my_rom(6022); 
 data6 <= my_rom(7377); 
 data7 <= my_rom(8732); 
 data8 <= my_rom(10087); 
 data9 <= my_rom(11442); 
 data10 <= my_rom(12797);
when "01001011011" => 
 data1 <= my_rom(603); 
 data2 <= my_rom(1958); 
 data3 <= my_rom(3313); 
 data4 <= my_rom(4668); 
 data5 <= my_rom(6023); 
 data6 <= my_rom(7378); 
 data7 <= my_rom(8733); 
 data8 <= my_rom(10088); 
 data9 <= my_rom(11443); 
 data10 <= my_rom(12798);
when "01001011100" => 
 data1 <= my_rom(604); 
 data2 <= my_rom(1959); 
 data3 <= my_rom(3314); 
 data4 <= my_rom(4669); 
 data5 <= my_rom(6024); 
 data6 <= my_rom(7379); 
 data7 <= my_rom(8734); 
 data8 <= my_rom(10089); 
 data9 <= my_rom(11444); 
 data10 <= my_rom(12799);
when "01001011101" => 
 data1 <= my_rom(605); 
 data2 <= my_rom(1960); 
 data3 <= my_rom(3315); 
 data4 <= my_rom(4670); 
 data5 <= my_rom(6025); 
 data6 <= my_rom(7380); 
 data7 <= my_rom(8735); 
 data8 <= my_rom(10090); 
 data9 <= my_rom(11445); 
 data10 <= my_rom(12800);
when "01001011110" => 
 data1 <= my_rom(606); 
 data2 <= my_rom(1961); 
 data3 <= my_rom(3316); 
 data4 <= my_rom(4671); 
 data5 <= my_rom(6026); 
 data6 <= my_rom(7381); 
 data7 <= my_rom(8736); 
 data8 <= my_rom(10091); 
 data9 <= my_rom(11446); 
 data10 <= my_rom(12801);
when "01001011111" => 
 data1 <= my_rom(607); 
 data2 <= my_rom(1962); 
 data3 <= my_rom(3317); 
 data4 <= my_rom(4672); 
 data5 <= my_rom(6027); 
 data6 <= my_rom(7382); 
 data7 <= my_rom(8737); 
 data8 <= my_rom(10092); 
 data9 <= my_rom(11447); 
 data10 <= my_rom(12802);
when "01001100000" => 
 data1 <= my_rom(608); 
 data2 <= my_rom(1963); 
 data3 <= my_rom(3318); 
 data4 <= my_rom(4673); 
 data5 <= my_rom(6028); 
 data6 <= my_rom(7383); 
 data7 <= my_rom(8738); 
 data8 <= my_rom(10093); 
 data9 <= my_rom(11448); 
 data10 <= my_rom(12803);
when "01001100001" => 
 data1 <= my_rom(609); 
 data2 <= my_rom(1964); 
 data3 <= my_rom(3319); 
 data4 <= my_rom(4674); 
 data5 <= my_rom(6029); 
 data6 <= my_rom(7384); 
 data7 <= my_rom(8739); 
 data8 <= my_rom(10094); 
 data9 <= my_rom(11449); 
 data10 <= my_rom(12804);
when "01001100010" => 
 data1 <= my_rom(610); 
 data2 <= my_rom(1965); 
 data3 <= my_rom(3320); 
 data4 <= my_rom(4675); 
 data5 <= my_rom(6030); 
 data6 <= my_rom(7385); 
 data7 <= my_rom(8740); 
 data8 <= my_rom(10095); 
 data9 <= my_rom(11450); 
 data10 <= my_rom(12805);
when "01001100011" => 
 data1 <= my_rom(611); 
 data2 <= my_rom(1966); 
 data3 <= my_rom(3321); 
 data4 <= my_rom(4676); 
 data5 <= my_rom(6031); 
 data6 <= my_rom(7386); 
 data7 <= my_rom(8741); 
 data8 <= my_rom(10096); 
 data9 <= my_rom(11451); 
 data10 <= my_rom(12806);
when "01001100100" => 
 data1 <= my_rom(612); 
 data2 <= my_rom(1967); 
 data3 <= my_rom(3322); 
 data4 <= my_rom(4677); 
 data5 <= my_rom(6032); 
 data6 <= my_rom(7387); 
 data7 <= my_rom(8742); 
 data8 <= my_rom(10097); 
 data9 <= my_rom(11452); 
 data10 <= my_rom(12807);
when "01001100101" => 
 data1 <= my_rom(613); 
 data2 <= my_rom(1968); 
 data3 <= my_rom(3323); 
 data4 <= my_rom(4678); 
 data5 <= my_rom(6033); 
 data6 <= my_rom(7388); 
 data7 <= my_rom(8743); 
 data8 <= my_rom(10098); 
 data9 <= my_rom(11453); 
 data10 <= my_rom(12808);
when "01001100110" => 
 data1 <= my_rom(614); 
 data2 <= my_rom(1969); 
 data3 <= my_rom(3324); 
 data4 <= my_rom(4679); 
 data5 <= my_rom(6034); 
 data6 <= my_rom(7389); 
 data7 <= my_rom(8744); 
 data8 <= my_rom(10099); 
 data9 <= my_rom(11454); 
 data10 <= my_rom(12809);
when "01001100111" => 
 data1 <= my_rom(615); 
 data2 <= my_rom(1970); 
 data3 <= my_rom(3325); 
 data4 <= my_rom(4680); 
 data5 <= my_rom(6035); 
 data6 <= my_rom(7390); 
 data7 <= my_rom(8745); 
 data8 <= my_rom(10100); 
 data9 <= my_rom(11455); 
 data10 <= my_rom(12810);
when "01001101000" => 
 data1 <= my_rom(616); 
 data2 <= my_rom(1971); 
 data3 <= my_rom(3326); 
 data4 <= my_rom(4681); 
 data5 <= my_rom(6036); 
 data6 <= my_rom(7391); 
 data7 <= my_rom(8746); 
 data8 <= my_rom(10101); 
 data9 <= my_rom(11456); 
 data10 <= my_rom(12811);
when "01001101001" => 
 data1 <= my_rom(617); 
 data2 <= my_rom(1972); 
 data3 <= my_rom(3327); 
 data4 <= my_rom(4682); 
 data5 <= my_rom(6037); 
 data6 <= my_rom(7392); 
 data7 <= my_rom(8747); 
 data8 <= my_rom(10102); 
 data9 <= my_rom(11457); 
 data10 <= my_rom(12812);
when "01001101010" => 
 data1 <= my_rom(618); 
 data2 <= my_rom(1973); 
 data3 <= my_rom(3328); 
 data4 <= my_rom(4683); 
 data5 <= my_rom(6038); 
 data6 <= my_rom(7393); 
 data7 <= my_rom(8748); 
 data8 <= my_rom(10103); 
 data9 <= my_rom(11458); 
 data10 <= my_rom(12813);
when "01001101011" => 
 data1 <= my_rom(619); 
 data2 <= my_rom(1974); 
 data3 <= my_rom(3329); 
 data4 <= my_rom(4684); 
 data5 <= my_rom(6039); 
 data6 <= my_rom(7394); 
 data7 <= my_rom(8749); 
 data8 <= my_rom(10104); 
 data9 <= my_rom(11459); 
 data10 <= my_rom(12814);
when "01001101100" => 
 data1 <= my_rom(620); 
 data2 <= my_rom(1975); 
 data3 <= my_rom(3330); 
 data4 <= my_rom(4685); 
 data5 <= my_rom(6040); 
 data6 <= my_rom(7395); 
 data7 <= my_rom(8750); 
 data8 <= my_rom(10105); 
 data9 <= my_rom(11460); 
 data10 <= my_rom(12815);
when "01001101101" => 
 data1 <= my_rom(621); 
 data2 <= my_rom(1976); 
 data3 <= my_rom(3331); 
 data4 <= my_rom(4686); 
 data5 <= my_rom(6041); 
 data6 <= my_rom(7396); 
 data7 <= my_rom(8751); 
 data8 <= my_rom(10106); 
 data9 <= my_rom(11461); 
 data10 <= my_rom(12816);
when "01001101110" => 
 data1 <= my_rom(622); 
 data2 <= my_rom(1977); 
 data3 <= my_rom(3332); 
 data4 <= my_rom(4687); 
 data5 <= my_rom(6042); 
 data6 <= my_rom(7397); 
 data7 <= my_rom(8752); 
 data8 <= my_rom(10107); 
 data9 <= my_rom(11462); 
 data10 <= my_rom(12817);
when "01001101111" => 
 data1 <= my_rom(623); 
 data2 <= my_rom(1978); 
 data3 <= my_rom(3333); 
 data4 <= my_rom(4688); 
 data5 <= my_rom(6043); 
 data6 <= my_rom(7398); 
 data7 <= my_rom(8753); 
 data8 <= my_rom(10108); 
 data9 <= my_rom(11463); 
 data10 <= my_rom(12818);
when "01001110000" => 
 data1 <= my_rom(624); 
 data2 <= my_rom(1979); 
 data3 <= my_rom(3334); 
 data4 <= my_rom(4689); 
 data5 <= my_rom(6044); 
 data6 <= my_rom(7399); 
 data7 <= my_rom(8754); 
 data8 <= my_rom(10109); 
 data9 <= my_rom(11464); 
 data10 <= my_rom(12819);
when "01001110001" => 
 data1 <= my_rom(625); 
 data2 <= my_rom(1980); 
 data3 <= my_rom(3335); 
 data4 <= my_rom(4690); 
 data5 <= my_rom(6045); 
 data6 <= my_rom(7400); 
 data7 <= my_rom(8755); 
 data8 <= my_rom(10110); 
 data9 <= my_rom(11465); 
 data10 <= my_rom(12820);
when "01001110010" => 
 data1 <= my_rom(626); 
 data2 <= my_rom(1981); 
 data3 <= my_rom(3336); 
 data4 <= my_rom(4691); 
 data5 <= my_rom(6046); 
 data6 <= my_rom(7401); 
 data7 <= my_rom(8756); 
 data8 <= my_rom(10111); 
 data9 <= my_rom(11466); 
 data10 <= my_rom(12821);
when "01001110011" => 
 data1 <= my_rom(627); 
 data2 <= my_rom(1982); 
 data3 <= my_rom(3337); 
 data4 <= my_rom(4692); 
 data5 <= my_rom(6047); 
 data6 <= my_rom(7402); 
 data7 <= my_rom(8757); 
 data8 <= my_rom(10112); 
 data9 <= my_rom(11467); 
 data10 <= my_rom(12822);
when "01001110100" => 
 data1 <= my_rom(628); 
 data2 <= my_rom(1983); 
 data3 <= my_rom(3338); 
 data4 <= my_rom(4693); 
 data5 <= my_rom(6048); 
 data6 <= my_rom(7403); 
 data7 <= my_rom(8758); 
 data8 <= my_rom(10113); 
 data9 <= my_rom(11468); 
 data10 <= my_rom(12823);
when "01001110101" => 
 data1 <= my_rom(629); 
 data2 <= my_rom(1984); 
 data3 <= my_rom(3339); 
 data4 <= my_rom(4694); 
 data5 <= my_rom(6049); 
 data6 <= my_rom(7404); 
 data7 <= my_rom(8759); 
 data8 <= my_rom(10114); 
 data9 <= my_rom(11469); 
 data10 <= my_rom(12824);
when "01001110110" => 
 data1 <= my_rom(630); 
 data2 <= my_rom(1985); 
 data3 <= my_rom(3340); 
 data4 <= my_rom(4695); 
 data5 <= my_rom(6050); 
 data6 <= my_rom(7405); 
 data7 <= my_rom(8760); 
 data8 <= my_rom(10115); 
 data9 <= my_rom(11470); 
 data10 <= my_rom(12825);
when "01001110111" => 
 data1 <= my_rom(631); 
 data2 <= my_rom(1986); 
 data3 <= my_rom(3341); 
 data4 <= my_rom(4696); 
 data5 <= my_rom(6051); 
 data6 <= my_rom(7406); 
 data7 <= my_rom(8761); 
 data8 <= my_rom(10116); 
 data9 <= my_rom(11471); 
 data10 <= my_rom(12826);
when "01001111000" => 
 data1 <= my_rom(632); 
 data2 <= my_rom(1987); 
 data3 <= my_rom(3342); 
 data4 <= my_rom(4697); 
 data5 <= my_rom(6052); 
 data6 <= my_rom(7407); 
 data7 <= my_rom(8762); 
 data8 <= my_rom(10117); 
 data9 <= my_rom(11472); 
 data10 <= my_rom(12827);
when "01001111001" => 
 data1 <= my_rom(633); 
 data2 <= my_rom(1988); 
 data3 <= my_rom(3343); 
 data4 <= my_rom(4698); 
 data5 <= my_rom(6053); 
 data6 <= my_rom(7408); 
 data7 <= my_rom(8763); 
 data8 <= my_rom(10118); 
 data9 <= my_rom(11473); 
 data10 <= my_rom(12828);
when "01001111010" => 
 data1 <= my_rom(634); 
 data2 <= my_rom(1989); 
 data3 <= my_rom(3344); 
 data4 <= my_rom(4699); 
 data5 <= my_rom(6054); 
 data6 <= my_rom(7409); 
 data7 <= my_rom(8764); 
 data8 <= my_rom(10119); 
 data9 <= my_rom(11474); 
 data10 <= my_rom(12829);
when "01001111011" => 
 data1 <= my_rom(635); 
 data2 <= my_rom(1990); 
 data3 <= my_rom(3345); 
 data4 <= my_rom(4700); 
 data5 <= my_rom(6055); 
 data6 <= my_rom(7410); 
 data7 <= my_rom(8765); 
 data8 <= my_rom(10120); 
 data9 <= my_rom(11475); 
 data10 <= my_rom(12830);
when "01001111100" => 
 data1 <= my_rom(636); 
 data2 <= my_rom(1991); 
 data3 <= my_rom(3346); 
 data4 <= my_rom(4701); 
 data5 <= my_rom(6056); 
 data6 <= my_rom(7411); 
 data7 <= my_rom(8766); 
 data8 <= my_rom(10121); 
 data9 <= my_rom(11476); 
 data10 <= my_rom(12831);
when "01001111101" => 
 data1 <= my_rom(637); 
 data2 <= my_rom(1992); 
 data3 <= my_rom(3347); 
 data4 <= my_rom(4702); 
 data5 <= my_rom(6057); 
 data6 <= my_rom(7412); 
 data7 <= my_rom(8767); 
 data8 <= my_rom(10122); 
 data9 <= my_rom(11477); 
 data10 <= my_rom(12832);
when "01001111110" => 
 data1 <= my_rom(638); 
 data2 <= my_rom(1993); 
 data3 <= my_rom(3348); 
 data4 <= my_rom(4703); 
 data5 <= my_rom(6058); 
 data6 <= my_rom(7413); 
 data7 <= my_rom(8768); 
 data8 <= my_rom(10123); 
 data9 <= my_rom(11478); 
 data10 <= my_rom(12833);
when "01001111111" => 
 data1 <= my_rom(639); 
 data2 <= my_rom(1994); 
 data3 <= my_rom(3349); 
 data4 <= my_rom(4704); 
 data5 <= my_rom(6059); 
 data6 <= my_rom(7414); 
 data7 <= my_rom(8769); 
 data8 <= my_rom(10124); 
 data9 <= my_rom(11479); 
 data10 <= my_rom(12834);
when "01010000000" => 
 data1 <= my_rom(640); 
 data2 <= my_rom(1995); 
 data3 <= my_rom(3350); 
 data4 <= my_rom(4705); 
 data5 <= my_rom(6060); 
 data6 <= my_rom(7415); 
 data7 <= my_rom(8770); 
 data8 <= my_rom(10125); 
 data9 <= my_rom(11480); 
 data10 <= my_rom(12835);
when "01010000001" => 
 data1 <= my_rom(641); 
 data2 <= my_rom(1996); 
 data3 <= my_rom(3351); 
 data4 <= my_rom(4706); 
 data5 <= my_rom(6061); 
 data6 <= my_rom(7416); 
 data7 <= my_rom(8771); 
 data8 <= my_rom(10126); 
 data9 <= my_rom(11481); 
 data10 <= my_rom(12836);
when "01010000010" => 
 data1 <= my_rom(642); 
 data2 <= my_rom(1997); 
 data3 <= my_rom(3352); 
 data4 <= my_rom(4707); 
 data5 <= my_rom(6062); 
 data6 <= my_rom(7417); 
 data7 <= my_rom(8772); 
 data8 <= my_rom(10127); 
 data9 <= my_rom(11482); 
 data10 <= my_rom(12837);
when "01010000011" => 
 data1 <= my_rom(643); 
 data2 <= my_rom(1998); 
 data3 <= my_rom(3353); 
 data4 <= my_rom(4708); 
 data5 <= my_rom(6063); 
 data6 <= my_rom(7418); 
 data7 <= my_rom(8773); 
 data8 <= my_rom(10128); 
 data9 <= my_rom(11483); 
 data10 <= my_rom(12838);
when "01010000100" => 
 data1 <= my_rom(644); 
 data2 <= my_rom(1999); 
 data3 <= my_rom(3354); 
 data4 <= my_rom(4709); 
 data5 <= my_rom(6064); 
 data6 <= my_rom(7419); 
 data7 <= my_rom(8774); 
 data8 <= my_rom(10129); 
 data9 <= my_rom(11484); 
 data10 <= my_rom(12839);
when "01010000101" => 
 data1 <= my_rom(645); 
 data2 <= my_rom(2000); 
 data3 <= my_rom(3355); 
 data4 <= my_rom(4710); 
 data5 <= my_rom(6065); 
 data6 <= my_rom(7420); 
 data7 <= my_rom(8775); 
 data8 <= my_rom(10130); 
 data9 <= my_rom(11485); 
 data10 <= my_rom(12840);
when "01010000110" => 
 data1 <= my_rom(646); 
 data2 <= my_rom(2001); 
 data3 <= my_rom(3356); 
 data4 <= my_rom(4711); 
 data5 <= my_rom(6066); 
 data6 <= my_rom(7421); 
 data7 <= my_rom(8776); 
 data8 <= my_rom(10131); 
 data9 <= my_rom(11486); 
 data10 <= my_rom(12841);
when "01010000111" => 
 data1 <= my_rom(647); 
 data2 <= my_rom(2002); 
 data3 <= my_rom(3357); 
 data4 <= my_rom(4712); 
 data5 <= my_rom(6067); 
 data6 <= my_rom(7422); 
 data7 <= my_rom(8777); 
 data8 <= my_rom(10132); 
 data9 <= my_rom(11487); 
 data10 <= my_rom(12842);
when "01010001000" => 
 data1 <= my_rom(648); 
 data2 <= my_rom(2003); 
 data3 <= my_rom(3358); 
 data4 <= my_rom(4713); 
 data5 <= my_rom(6068); 
 data6 <= my_rom(7423); 
 data7 <= my_rom(8778); 
 data8 <= my_rom(10133); 
 data9 <= my_rom(11488); 
 data10 <= my_rom(12843);
when "01010001001" => 
 data1 <= my_rom(649); 
 data2 <= my_rom(2004); 
 data3 <= my_rom(3359); 
 data4 <= my_rom(4714); 
 data5 <= my_rom(6069); 
 data6 <= my_rom(7424); 
 data7 <= my_rom(8779); 
 data8 <= my_rom(10134); 
 data9 <= my_rom(11489); 
 data10 <= my_rom(12844);
when "01010001010" => 
 data1 <= my_rom(650); 
 data2 <= my_rom(2005); 
 data3 <= my_rom(3360); 
 data4 <= my_rom(4715); 
 data5 <= my_rom(6070); 
 data6 <= my_rom(7425); 
 data7 <= my_rom(8780); 
 data8 <= my_rom(10135); 
 data9 <= my_rom(11490); 
 data10 <= my_rom(12845);
when "01010001011" => 
 data1 <= my_rom(651); 
 data2 <= my_rom(2006); 
 data3 <= my_rom(3361); 
 data4 <= my_rom(4716); 
 data5 <= my_rom(6071); 
 data6 <= my_rom(7426); 
 data7 <= my_rom(8781); 
 data8 <= my_rom(10136); 
 data9 <= my_rom(11491); 
 data10 <= my_rom(12846);
when "01010001100" => 
 data1 <= my_rom(652); 
 data2 <= my_rom(2007); 
 data3 <= my_rom(3362); 
 data4 <= my_rom(4717); 
 data5 <= my_rom(6072); 
 data6 <= my_rom(7427); 
 data7 <= my_rom(8782); 
 data8 <= my_rom(10137); 
 data9 <= my_rom(11492); 
 data10 <= my_rom(12847);
when "01010001101" => 
 data1 <= my_rom(653); 
 data2 <= my_rom(2008); 
 data3 <= my_rom(3363); 
 data4 <= my_rom(4718); 
 data5 <= my_rom(6073); 
 data6 <= my_rom(7428); 
 data7 <= my_rom(8783); 
 data8 <= my_rom(10138); 
 data9 <= my_rom(11493); 
 data10 <= my_rom(12848);
when "01010001110" => 
 data1 <= my_rom(654); 
 data2 <= my_rom(2009); 
 data3 <= my_rom(3364); 
 data4 <= my_rom(4719); 
 data5 <= my_rom(6074); 
 data6 <= my_rom(7429); 
 data7 <= my_rom(8784); 
 data8 <= my_rom(10139); 
 data9 <= my_rom(11494); 
 data10 <= my_rom(12849);
when "01010001111" => 
 data1 <= my_rom(655); 
 data2 <= my_rom(2010); 
 data3 <= my_rom(3365); 
 data4 <= my_rom(4720); 
 data5 <= my_rom(6075); 
 data6 <= my_rom(7430); 
 data7 <= my_rom(8785); 
 data8 <= my_rom(10140); 
 data9 <= my_rom(11495); 
 data10 <= my_rom(12850);
when "01010010000" => 
 data1 <= my_rom(656); 
 data2 <= my_rom(2011); 
 data3 <= my_rom(3366); 
 data4 <= my_rom(4721); 
 data5 <= my_rom(6076); 
 data6 <= my_rom(7431); 
 data7 <= my_rom(8786); 
 data8 <= my_rom(10141); 
 data9 <= my_rom(11496); 
 data10 <= my_rom(12851);
when "01010010001" => 
 data1 <= my_rom(657); 
 data2 <= my_rom(2012); 
 data3 <= my_rom(3367); 
 data4 <= my_rom(4722); 
 data5 <= my_rom(6077); 
 data6 <= my_rom(7432); 
 data7 <= my_rom(8787); 
 data8 <= my_rom(10142); 
 data9 <= my_rom(11497); 
 data10 <= my_rom(12852);
when "01010010010" => 
 data1 <= my_rom(658); 
 data2 <= my_rom(2013); 
 data3 <= my_rom(3368); 
 data4 <= my_rom(4723); 
 data5 <= my_rom(6078); 
 data6 <= my_rom(7433); 
 data7 <= my_rom(8788); 
 data8 <= my_rom(10143); 
 data9 <= my_rom(11498); 
 data10 <= my_rom(12853);
when "01010010011" => 
 data1 <= my_rom(659); 
 data2 <= my_rom(2014); 
 data3 <= my_rom(3369); 
 data4 <= my_rom(4724); 
 data5 <= my_rom(6079); 
 data6 <= my_rom(7434); 
 data7 <= my_rom(8789); 
 data8 <= my_rom(10144); 
 data9 <= my_rom(11499); 
 data10 <= my_rom(12854);
when "01010010100" => 
 data1 <= my_rom(660); 
 data2 <= my_rom(2015); 
 data3 <= my_rom(3370); 
 data4 <= my_rom(4725); 
 data5 <= my_rom(6080); 
 data6 <= my_rom(7435); 
 data7 <= my_rom(8790); 
 data8 <= my_rom(10145); 
 data9 <= my_rom(11500); 
 data10 <= my_rom(12855);
when "01010010101" => 
 data1 <= my_rom(661); 
 data2 <= my_rom(2016); 
 data3 <= my_rom(3371); 
 data4 <= my_rom(4726); 
 data5 <= my_rom(6081); 
 data6 <= my_rom(7436); 
 data7 <= my_rom(8791); 
 data8 <= my_rom(10146); 
 data9 <= my_rom(11501); 
 data10 <= my_rom(12856);
when "01010010110" => 
 data1 <= my_rom(662); 
 data2 <= my_rom(2017); 
 data3 <= my_rom(3372); 
 data4 <= my_rom(4727); 
 data5 <= my_rom(6082); 
 data6 <= my_rom(7437); 
 data7 <= my_rom(8792); 
 data8 <= my_rom(10147); 
 data9 <= my_rom(11502); 
 data10 <= my_rom(12857);
when "01010010111" => 
 data1 <= my_rom(663); 
 data2 <= my_rom(2018); 
 data3 <= my_rom(3373); 
 data4 <= my_rom(4728); 
 data5 <= my_rom(6083); 
 data6 <= my_rom(7438); 
 data7 <= my_rom(8793); 
 data8 <= my_rom(10148); 
 data9 <= my_rom(11503); 
 data10 <= my_rom(12858);
when "01010011000" => 
 data1 <= my_rom(664); 
 data2 <= my_rom(2019); 
 data3 <= my_rom(3374); 
 data4 <= my_rom(4729); 
 data5 <= my_rom(6084); 
 data6 <= my_rom(7439); 
 data7 <= my_rom(8794); 
 data8 <= my_rom(10149); 
 data9 <= my_rom(11504); 
 data10 <= my_rom(12859);
when "01010011001" => 
 data1 <= my_rom(665); 
 data2 <= my_rom(2020); 
 data3 <= my_rom(3375); 
 data4 <= my_rom(4730); 
 data5 <= my_rom(6085); 
 data6 <= my_rom(7440); 
 data7 <= my_rom(8795); 
 data8 <= my_rom(10150); 
 data9 <= my_rom(11505); 
 data10 <= my_rom(12860);
when "01010011010" => 
 data1 <= my_rom(666); 
 data2 <= my_rom(2021); 
 data3 <= my_rom(3376); 
 data4 <= my_rom(4731); 
 data5 <= my_rom(6086); 
 data6 <= my_rom(7441); 
 data7 <= my_rom(8796); 
 data8 <= my_rom(10151); 
 data9 <= my_rom(11506); 
 data10 <= my_rom(12861);
when "01010011011" => 
 data1 <= my_rom(667); 
 data2 <= my_rom(2022); 
 data3 <= my_rom(3377); 
 data4 <= my_rom(4732); 
 data5 <= my_rom(6087); 
 data6 <= my_rom(7442); 
 data7 <= my_rom(8797); 
 data8 <= my_rom(10152); 
 data9 <= my_rom(11507); 
 data10 <= my_rom(12862);
when "01010011100" => 
 data1 <= my_rom(668); 
 data2 <= my_rom(2023); 
 data3 <= my_rom(3378); 
 data4 <= my_rom(4733); 
 data5 <= my_rom(6088); 
 data6 <= my_rom(7443); 
 data7 <= my_rom(8798); 
 data8 <= my_rom(10153); 
 data9 <= my_rom(11508); 
 data10 <= my_rom(12863);
when "01010011101" => 
 data1 <= my_rom(669); 
 data2 <= my_rom(2024); 
 data3 <= my_rom(3379); 
 data4 <= my_rom(4734); 
 data5 <= my_rom(6089); 
 data6 <= my_rom(7444); 
 data7 <= my_rom(8799); 
 data8 <= my_rom(10154); 
 data9 <= my_rom(11509); 
 data10 <= my_rom(12864);
when "01010011110" => 
 data1 <= my_rom(670); 
 data2 <= my_rom(2025); 
 data3 <= my_rom(3380); 
 data4 <= my_rom(4735); 
 data5 <= my_rom(6090); 
 data6 <= my_rom(7445); 
 data7 <= my_rom(8800); 
 data8 <= my_rom(10155); 
 data9 <= my_rom(11510); 
 data10 <= my_rom(12865);
when "01010011111" => 
 data1 <= my_rom(671); 
 data2 <= my_rom(2026); 
 data3 <= my_rom(3381); 
 data4 <= my_rom(4736); 
 data5 <= my_rom(6091); 
 data6 <= my_rom(7446); 
 data7 <= my_rom(8801); 
 data8 <= my_rom(10156); 
 data9 <= my_rom(11511); 
 data10 <= my_rom(12866);
when "01010100000" => 
 data1 <= my_rom(672); 
 data2 <= my_rom(2027); 
 data3 <= my_rom(3382); 
 data4 <= my_rom(4737); 
 data5 <= my_rom(6092); 
 data6 <= my_rom(7447); 
 data7 <= my_rom(8802); 
 data8 <= my_rom(10157); 
 data9 <= my_rom(11512); 
 data10 <= my_rom(12867);
when "01010100001" => 
 data1 <= my_rom(673); 
 data2 <= my_rom(2028); 
 data3 <= my_rom(3383); 
 data4 <= my_rom(4738); 
 data5 <= my_rom(6093); 
 data6 <= my_rom(7448); 
 data7 <= my_rom(8803); 
 data8 <= my_rom(10158); 
 data9 <= my_rom(11513); 
 data10 <= my_rom(12868);
when "01010100010" => 
 data1 <= my_rom(674); 
 data2 <= my_rom(2029); 
 data3 <= my_rom(3384); 
 data4 <= my_rom(4739); 
 data5 <= my_rom(6094); 
 data6 <= my_rom(7449); 
 data7 <= my_rom(8804); 
 data8 <= my_rom(10159); 
 data9 <= my_rom(11514); 
 data10 <= my_rom(12869);
when "01010100011" => 
 data1 <= my_rom(675); 
 data2 <= my_rom(2030); 
 data3 <= my_rom(3385); 
 data4 <= my_rom(4740); 
 data5 <= my_rom(6095); 
 data6 <= my_rom(7450); 
 data7 <= my_rom(8805); 
 data8 <= my_rom(10160); 
 data9 <= my_rom(11515); 
 data10 <= my_rom(12870);
when "01010100100" => 
 data1 <= my_rom(676); 
 data2 <= my_rom(2031); 
 data3 <= my_rom(3386); 
 data4 <= my_rom(4741); 
 data5 <= my_rom(6096); 
 data6 <= my_rom(7451); 
 data7 <= my_rom(8806); 
 data8 <= my_rom(10161); 
 data9 <= my_rom(11516); 
 data10 <= my_rom(12871);
when "01010100101" => 
 data1 <= my_rom(677); 
 data2 <= my_rom(2032); 
 data3 <= my_rom(3387); 
 data4 <= my_rom(4742); 
 data5 <= my_rom(6097); 
 data6 <= my_rom(7452); 
 data7 <= my_rom(8807); 
 data8 <= my_rom(10162); 
 data9 <= my_rom(11517); 
 data10 <= my_rom(12872);
when "01010100110" => 
 data1 <= my_rom(678); 
 data2 <= my_rom(2033); 
 data3 <= my_rom(3388); 
 data4 <= my_rom(4743); 
 data5 <= my_rom(6098); 
 data6 <= my_rom(7453); 
 data7 <= my_rom(8808); 
 data8 <= my_rom(10163); 
 data9 <= my_rom(11518); 
 data10 <= my_rom(12873);
when "01010100111" => 
 data1 <= my_rom(679); 
 data2 <= my_rom(2034); 
 data3 <= my_rom(3389); 
 data4 <= my_rom(4744); 
 data5 <= my_rom(6099); 
 data6 <= my_rom(7454); 
 data7 <= my_rom(8809); 
 data8 <= my_rom(10164); 
 data9 <= my_rom(11519); 
 data10 <= my_rom(12874);
when "01010101000" => 
 data1 <= my_rom(680); 
 data2 <= my_rom(2035); 
 data3 <= my_rom(3390); 
 data4 <= my_rom(4745); 
 data5 <= my_rom(6100); 
 data6 <= my_rom(7455); 
 data7 <= my_rom(8810); 
 data8 <= my_rom(10165); 
 data9 <= my_rom(11520); 
 data10 <= my_rom(12875);
when "01010101001" => 
 data1 <= my_rom(681); 
 data2 <= my_rom(2036); 
 data3 <= my_rom(3391); 
 data4 <= my_rom(4746); 
 data5 <= my_rom(6101); 
 data6 <= my_rom(7456); 
 data7 <= my_rom(8811); 
 data8 <= my_rom(10166); 
 data9 <= my_rom(11521); 
 data10 <= my_rom(12876);
when "01010101010" => 
 data1 <= my_rom(682); 
 data2 <= my_rom(2037); 
 data3 <= my_rom(3392); 
 data4 <= my_rom(4747); 
 data5 <= my_rom(6102); 
 data6 <= my_rom(7457); 
 data7 <= my_rom(8812); 
 data8 <= my_rom(10167); 
 data9 <= my_rom(11522); 
 data10 <= my_rom(12877);
when "01010101011" => 
 data1 <= my_rom(683); 
 data2 <= my_rom(2038); 
 data3 <= my_rom(3393); 
 data4 <= my_rom(4748); 
 data5 <= my_rom(6103); 
 data6 <= my_rom(7458); 
 data7 <= my_rom(8813); 
 data8 <= my_rom(10168); 
 data9 <= my_rom(11523); 
 data10 <= my_rom(12878);
when "01010101100" => 
 data1 <= my_rom(684); 
 data2 <= my_rom(2039); 
 data3 <= my_rom(3394); 
 data4 <= my_rom(4749); 
 data5 <= my_rom(6104); 
 data6 <= my_rom(7459); 
 data7 <= my_rom(8814); 
 data8 <= my_rom(10169); 
 data9 <= my_rom(11524); 
 data10 <= my_rom(12879);
when "01010101101" => 
 data1 <= my_rom(685); 
 data2 <= my_rom(2040); 
 data3 <= my_rom(3395); 
 data4 <= my_rom(4750); 
 data5 <= my_rom(6105); 
 data6 <= my_rom(7460); 
 data7 <= my_rom(8815); 
 data8 <= my_rom(10170); 
 data9 <= my_rom(11525); 
 data10 <= my_rom(12880);
when "01010101110" => 
 data1 <= my_rom(686); 
 data2 <= my_rom(2041); 
 data3 <= my_rom(3396); 
 data4 <= my_rom(4751); 
 data5 <= my_rom(6106); 
 data6 <= my_rom(7461); 
 data7 <= my_rom(8816); 
 data8 <= my_rom(10171); 
 data9 <= my_rom(11526); 
 data10 <= my_rom(12881);
when "01010101111" => 
 data1 <= my_rom(687); 
 data2 <= my_rom(2042); 
 data3 <= my_rom(3397); 
 data4 <= my_rom(4752); 
 data5 <= my_rom(6107); 
 data6 <= my_rom(7462); 
 data7 <= my_rom(8817); 
 data8 <= my_rom(10172); 
 data9 <= my_rom(11527); 
 data10 <= my_rom(12882);
when "01010110000" => 
 data1 <= my_rom(688); 
 data2 <= my_rom(2043); 
 data3 <= my_rom(3398); 
 data4 <= my_rom(4753); 
 data5 <= my_rom(6108); 
 data6 <= my_rom(7463); 
 data7 <= my_rom(8818); 
 data8 <= my_rom(10173); 
 data9 <= my_rom(11528); 
 data10 <= my_rom(12883);
when "01010110001" => 
 data1 <= my_rom(689); 
 data2 <= my_rom(2044); 
 data3 <= my_rom(3399); 
 data4 <= my_rom(4754); 
 data5 <= my_rom(6109); 
 data6 <= my_rom(7464); 
 data7 <= my_rom(8819); 
 data8 <= my_rom(10174); 
 data9 <= my_rom(11529); 
 data10 <= my_rom(12884);
when "01010110010" => 
 data1 <= my_rom(690); 
 data2 <= my_rom(2045); 
 data3 <= my_rom(3400); 
 data4 <= my_rom(4755); 
 data5 <= my_rom(6110); 
 data6 <= my_rom(7465); 
 data7 <= my_rom(8820); 
 data8 <= my_rom(10175); 
 data9 <= my_rom(11530); 
 data10 <= my_rom(12885);
when "01010110011" => 
 data1 <= my_rom(691); 
 data2 <= my_rom(2046); 
 data3 <= my_rom(3401); 
 data4 <= my_rom(4756); 
 data5 <= my_rom(6111); 
 data6 <= my_rom(7466); 
 data7 <= my_rom(8821); 
 data8 <= my_rom(10176); 
 data9 <= my_rom(11531); 
 data10 <= my_rom(12886);
when "01010110100" => 
 data1 <= my_rom(692); 
 data2 <= my_rom(2047); 
 data3 <= my_rom(3402); 
 data4 <= my_rom(4757); 
 data5 <= my_rom(6112); 
 data6 <= my_rom(7467); 
 data7 <= my_rom(8822); 
 data8 <= my_rom(10177); 
 data9 <= my_rom(11532); 
 data10 <= my_rom(12887);
when "01010110101" => 
 data1 <= my_rom(693); 
 data2 <= my_rom(2048); 
 data3 <= my_rom(3403); 
 data4 <= my_rom(4758); 
 data5 <= my_rom(6113); 
 data6 <= my_rom(7468); 
 data7 <= my_rom(8823); 
 data8 <= my_rom(10178); 
 data9 <= my_rom(11533); 
 data10 <= my_rom(12888);
when "01010110110" => 
 data1 <= my_rom(694); 
 data2 <= my_rom(2049); 
 data3 <= my_rom(3404); 
 data4 <= my_rom(4759); 
 data5 <= my_rom(6114); 
 data6 <= my_rom(7469); 
 data7 <= my_rom(8824); 
 data8 <= my_rom(10179); 
 data9 <= my_rom(11534); 
 data10 <= my_rom(12889);
when "01010110111" => 
 data1 <= my_rom(695); 
 data2 <= my_rom(2050); 
 data3 <= my_rom(3405); 
 data4 <= my_rom(4760); 
 data5 <= my_rom(6115); 
 data6 <= my_rom(7470); 
 data7 <= my_rom(8825); 
 data8 <= my_rom(10180); 
 data9 <= my_rom(11535); 
 data10 <= my_rom(12890);
when "01010111000" => 
 data1 <= my_rom(696); 
 data2 <= my_rom(2051); 
 data3 <= my_rom(3406); 
 data4 <= my_rom(4761); 
 data5 <= my_rom(6116); 
 data6 <= my_rom(7471); 
 data7 <= my_rom(8826); 
 data8 <= my_rom(10181); 
 data9 <= my_rom(11536); 
 data10 <= my_rom(12891);
when "01010111001" => 
 data1 <= my_rom(697); 
 data2 <= my_rom(2052); 
 data3 <= my_rom(3407); 
 data4 <= my_rom(4762); 
 data5 <= my_rom(6117); 
 data6 <= my_rom(7472); 
 data7 <= my_rom(8827); 
 data8 <= my_rom(10182); 
 data9 <= my_rom(11537); 
 data10 <= my_rom(12892);
when "01010111010" => 
 data1 <= my_rom(698); 
 data2 <= my_rom(2053); 
 data3 <= my_rom(3408); 
 data4 <= my_rom(4763); 
 data5 <= my_rom(6118); 
 data6 <= my_rom(7473); 
 data7 <= my_rom(8828); 
 data8 <= my_rom(10183); 
 data9 <= my_rom(11538); 
 data10 <= my_rom(12893);
when "01010111011" => 
 data1 <= my_rom(699); 
 data2 <= my_rom(2054); 
 data3 <= my_rom(3409); 
 data4 <= my_rom(4764); 
 data5 <= my_rom(6119); 
 data6 <= my_rom(7474); 
 data7 <= my_rom(8829); 
 data8 <= my_rom(10184); 
 data9 <= my_rom(11539); 
 data10 <= my_rom(12894);
when "01010111100" => 
 data1 <= my_rom(700); 
 data2 <= my_rom(2055); 
 data3 <= my_rom(3410); 
 data4 <= my_rom(4765); 
 data5 <= my_rom(6120); 
 data6 <= my_rom(7475); 
 data7 <= my_rom(8830); 
 data8 <= my_rom(10185); 
 data9 <= my_rom(11540); 
 data10 <= my_rom(12895);
when "01010111101" => 
 data1 <= my_rom(701); 
 data2 <= my_rom(2056); 
 data3 <= my_rom(3411); 
 data4 <= my_rom(4766); 
 data5 <= my_rom(6121); 
 data6 <= my_rom(7476); 
 data7 <= my_rom(8831); 
 data8 <= my_rom(10186); 
 data9 <= my_rom(11541); 
 data10 <= my_rom(12896);
when "01010111110" => 
 data1 <= my_rom(702); 
 data2 <= my_rom(2057); 
 data3 <= my_rom(3412); 
 data4 <= my_rom(4767); 
 data5 <= my_rom(6122); 
 data6 <= my_rom(7477); 
 data7 <= my_rom(8832); 
 data8 <= my_rom(10187); 
 data9 <= my_rom(11542); 
 data10 <= my_rom(12897);
when "01010111111" => 
 data1 <= my_rom(703); 
 data2 <= my_rom(2058); 
 data3 <= my_rom(3413); 
 data4 <= my_rom(4768); 
 data5 <= my_rom(6123); 
 data6 <= my_rom(7478); 
 data7 <= my_rom(8833); 
 data8 <= my_rom(10188); 
 data9 <= my_rom(11543); 
 data10 <= my_rom(12898);
when "01011000000" => 
 data1 <= my_rom(704); 
 data2 <= my_rom(2059); 
 data3 <= my_rom(3414); 
 data4 <= my_rom(4769); 
 data5 <= my_rom(6124); 
 data6 <= my_rom(7479); 
 data7 <= my_rom(8834); 
 data8 <= my_rom(10189); 
 data9 <= my_rom(11544); 
 data10 <= my_rom(12899);
when "01011000001" => 
 data1 <= my_rom(705); 
 data2 <= my_rom(2060); 
 data3 <= my_rom(3415); 
 data4 <= my_rom(4770); 
 data5 <= my_rom(6125); 
 data6 <= my_rom(7480); 
 data7 <= my_rom(8835); 
 data8 <= my_rom(10190); 
 data9 <= my_rom(11545); 
 data10 <= my_rom(12900);
when "01011000010" => 
 data1 <= my_rom(706); 
 data2 <= my_rom(2061); 
 data3 <= my_rom(3416); 
 data4 <= my_rom(4771); 
 data5 <= my_rom(6126); 
 data6 <= my_rom(7481); 
 data7 <= my_rom(8836); 
 data8 <= my_rom(10191); 
 data9 <= my_rom(11546); 
 data10 <= my_rom(12901);
when "01011000011" => 
 data1 <= my_rom(707); 
 data2 <= my_rom(2062); 
 data3 <= my_rom(3417); 
 data4 <= my_rom(4772); 
 data5 <= my_rom(6127); 
 data6 <= my_rom(7482); 
 data7 <= my_rom(8837); 
 data8 <= my_rom(10192); 
 data9 <= my_rom(11547); 
 data10 <= my_rom(12902);
when "01011000100" => 
 data1 <= my_rom(708); 
 data2 <= my_rom(2063); 
 data3 <= my_rom(3418); 
 data4 <= my_rom(4773); 
 data5 <= my_rom(6128); 
 data6 <= my_rom(7483); 
 data7 <= my_rom(8838); 
 data8 <= my_rom(10193); 
 data9 <= my_rom(11548); 
 data10 <= my_rom(12903);
when "01011000101" => 
 data1 <= my_rom(709); 
 data2 <= my_rom(2064); 
 data3 <= my_rom(3419); 
 data4 <= my_rom(4774); 
 data5 <= my_rom(6129); 
 data6 <= my_rom(7484); 
 data7 <= my_rom(8839); 
 data8 <= my_rom(10194); 
 data9 <= my_rom(11549); 
 data10 <= my_rom(12904);
when "01011000110" => 
 data1 <= my_rom(710); 
 data2 <= my_rom(2065); 
 data3 <= my_rom(3420); 
 data4 <= my_rom(4775); 
 data5 <= my_rom(6130); 
 data6 <= my_rom(7485); 
 data7 <= my_rom(8840); 
 data8 <= my_rom(10195); 
 data9 <= my_rom(11550); 
 data10 <= my_rom(12905);
when "01011000111" => 
 data1 <= my_rom(711); 
 data2 <= my_rom(2066); 
 data3 <= my_rom(3421); 
 data4 <= my_rom(4776); 
 data5 <= my_rom(6131); 
 data6 <= my_rom(7486); 
 data7 <= my_rom(8841); 
 data8 <= my_rom(10196); 
 data9 <= my_rom(11551); 
 data10 <= my_rom(12906);
when "01011001000" => 
 data1 <= my_rom(712); 
 data2 <= my_rom(2067); 
 data3 <= my_rom(3422); 
 data4 <= my_rom(4777); 
 data5 <= my_rom(6132); 
 data6 <= my_rom(7487); 
 data7 <= my_rom(8842); 
 data8 <= my_rom(10197); 
 data9 <= my_rom(11552); 
 data10 <= my_rom(12907);
when "01011001001" => 
 data1 <= my_rom(713); 
 data2 <= my_rom(2068); 
 data3 <= my_rom(3423); 
 data4 <= my_rom(4778); 
 data5 <= my_rom(6133); 
 data6 <= my_rom(7488); 
 data7 <= my_rom(8843); 
 data8 <= my_rom(10198); 
 data9 <= my_rom(11553); 
 data10 <= my_rom(12908);
when "01011001010" => 
 data1 <= my_rom(714); 
 data2 <= my_rom(2069); 
 data3 <= my_rom(3424); 
 data4 <= my_rom(4779); 
 data5 <= my_rom(6134); 
 data6 <= my_rom(7489); 
 data7 <= my_rom(8844); 
 data8 <= my_rom(10199); 
 data9 <= my_rom(11554); 
 data10 <= my_rom(12909);
when "01011001011" => 
 data1 <= my_rom(715); 
 data2 <= my_rom(2070); 
 data3 <= my_rom(3425); 
 data4 <= my_rom(4780); 
 data5 <= my_rom(6135); 
 data6 <= my_rom(7490); 
 data7 <= my_rom(8845); 
 data8 <= my_rom(10200); 
 data9 <= my_rom(11555); 
 data10 <= my_rom(12910);
when "01011001100" => 
 data1 <= my_rom(716); 
 data2 <= my_rom(2071); 
 data3 <= my_rom(3426); 
 data4 <= my_rom(4781); 
 data5 <= my_rom(6136); 
 data6 <= my_rom(7491); 
 data7 <= my_rom(8846); 
 data8 <= my_rom(10201); 
 data9 <= my_rom(11556); 
 data10 <= my_rom(12911);
when "01011001101" => 
 data1 <= my_rom(717); 
 data2 <= my_rom(2072); 
 data3 <= my_rom(3427); 
 data4 <= my_rom(4782); 
 data5 <= my_rom(6137); 
 data6 <= my_rom(7492); 
 data7 <= my_rom(8847); 
 data8 <= my_rom(10202); 
 data9 <= my_rom(11557); 
 data10 <= my_rom(12912);
when "01011001110" => 
 data1 <= my_rom(718); 
 data2 <= my_rom(2073); 
 data3 <= my_rom(3428); 
 data4 <= my_rom(4783); 
 data5 <= my_rom(6138); 
 data6 <= my_rom(7493); 
 data7 <= my_rom(8848); 
 data8 <= my_rom(10203); 
 data9 <= my_rom(11558); 
 data10 <= my_rom(12913);
when "01011001111" => 
 data1 <= my_rom(719); 
 data2 <= my_rom(2074); 
 data3 <= my_rom(3429); 
 data4 <= my_rom(4784); 
 data5 <= my_rom(6139); 
 data6 <= my_rom(7494); 
 data7 <= my_rom(8849); 
 data8 <= my_rom(10204); 
 data9 <= my_rom(11559); 
 data10 <= my_rom(12914);
when "01011010000" => 
 data1 <= my_rom(720); 
 data2 <= my_rom(2075); 
 data3 <= my_rom(3430); 
 data4 <= my_rom(4785); 
 data5 <= my_rom(6140); 
 data6 <= my_rom(7495); 
 data7 <= my_rom(8850); 
 data8 <= my_rom(10205); 
 data9 <= my_rom(11560); 
 data10 <= my_rom(12915);
when "01011010001" => 
 data1 <= my_rom(721); 
 data2 <= my_rom(2076); 
 data3 <= my_rom(3431); 
 data4 <= my_rom(4786); 
 data5 <= my_rom(6141); 
 data6 <= my_rom(7496); 
 data7 <= my_rom(8851); 
 data8 <= my_rom(10206); 
 data9 <= my_rom(11561); 
 data10 <= my_rom(12916);
when "01011010010" => 
 data1 <= my_rom(722); 
 data2 <= my_rom(2077); 
 data3 <= my_rom(3432); 
 data4 <= my_rom(4787); 
 data5 <= my_rom(6142); 
 data6 <= my_rom(7497); 
 data7 <= my_rom(8852); 
 data8 <= my_rom(10207); 
 data9 <= my_rom(11562); 
 data10 <= my_rom(12917);
when "01011010011" => 
 data1 <= my_rom(723); 
 data2 <= my_rom(2078); 
 data3 <= my_rom(3433); 
 data4 <= my_rom(4788); 
 data5 <= my_rom(6143); 
 data6 <= my_rom(7498); 
 data7 <= my_rom(8853); 
 data8 <= my_rom(10208); 
 data9 <= my_rom(11563); 
 data10 <= my_rom(12918);
when "01011010100" => 
 data1 <= my_rom(724); 
 data2 <= my_rom(2079); 
 data3 <= my_rom(3434); 
 data4 <= my_rom(4789); 
 data5 <= my_rom(6144); 
 data6 <= my_rom(7499); 
 data7 <= my_rom(8854); 
 data8 <= my_rom(10209); 
 data9 <= my_rom(11564); 
 data10 <= my_rom(12919);
when "01011010101" => 
 data1 <= my_rom(725); 
 data2 <= my_rom(2080); 
 data3 <= my_rom(3435); 
 data4 <= my_rom(4790); 
 data5 <= my_rom(6145); 
 data6 <= my_rom(7500); 
 data7 <= my_rom(8855); 
 data8 <= my_rom(10210); 
 data9 <= my_rom(11565); 
 data10 <= my_rom(12920);
when "01011010110" => 
 data1 <= my_rom(726); 
 data2 <= my_rom(2081); 
 data3 <= my_rom(3436); 
 data4 <= my_rom(4791); 
 data5 <= my_rom(6146); 
 data6 <= my_rom(7501); 
 data7 <= my_rom(8856); 
 data8 <= my_rom(10211); 
 data9 <= my_rom(11566); 
 data10 <= my_rom(12921);
when "01011010111" => 
 data1 <= my_rom(727); 
 data2 <= my_rom(2082); 
 data3 <= my_rom(3437); 
 data4 <= my_rom(4792); 
 data5 <= my_rom(6147); 
 data6 <= my_rom(7502); 
 data7 <= my_rom(8857); 
 data8 <= my_rom(10212); 
 data9 <= my_rom(11567); 
 data10 <= my_rom(12922);
when "01011011000" => 
 data1 <= my_rom(728); 
 data2 <= my_rom(2083); 
 data3 <= my_rom(3438); 
 data4 <= my_rom(4793); 
 data5 <= my_rom(6148); 
 data6 <= my_rom(7503); 
 data7 <= my_rom(8858); 
 data8 <= my_rom(10213); 
 data9 <= my_rom(11568); 
 data10 <= my_rom(12923);
when "01011011001" => 
 data1 <= my_rom(729); 
 data2 <= my_rom(2084); 
 data3 <= my_rom(3439); 
 data4 <= my_rom(4794); 
 data5 <= my_rom(6149); 
 data6 <= my_rom(7504); 
 data7 <= my_rom(8859); 
 data8 <= my_rom(10214); 
 data9 <= my_rom(11569); 
 data10 <= my_rom(12924);
when "01011011010" => 
 data1 <= my_rom(730); 
 data2 <= my_rom(2085); 
 data3 <= my_rom(3440); 
 data4 <= my_rom(4795); 
 data5 <= my_rom(6150); 
 data6 <= my_rom(7505); 
 data7 <= my_rom(8860); 
 data8 <= my_rom(10215); 
 data9 <= my_rom(11570); 
 data10 <= my_rom(12925);
when "01011011011" => 
 data1 <= my_rom(731); 
 data2 <= my_rom(2086); 
 data3 <= my_rom(3441); 
 data4 <= my_rom(4796); 
 data5 <= my_rom(6151); 
 data6 <= my_rom(7506); 
 data7 <= my_rom(8861); 
 data8 <= my_rom(10216); 
 data9 <= my_rom(11571); 
 data10 <= my_rom(12926);
when "01011011100" => 
 data1 <= my_rom(732); 
 data2 <= my_rom(2087); 
 data3 <= my_rom(3442); 
 data4 <= my_rom(4797); 
 data5 <= my_rom(6152); 
 data6 <= my_rom(7507); 
 data7 <= my_rom(8862); 
 data8 <= my_rom(10217); 
 data9 <= my_rom(11572); 
 data10 <= my_rom(12927);
when "01011011101" => 
 data1 <= my_rom(733); 
 data2 <= my_rom(2088); 
 data3 <= my_rom(3443); 
 data4 <= my_rom(4798); 
 data5 <= my_rom(6153); 
 data6 <= my_rom(7508); 
 data7 <= my_rom(8863); 
 data8 <= my_rom(10218); 
 data9 <= my_rom(11573); 
 data10 <= my_rom(12928);
when "01011011110" => 
 data1 <= my_rom(734); 
 data2 <= my_rom(2089); 
 data3 <= my_rom(3444); 
 data4 <= my_rom(4799); 
 data5 <= my_rom(6154); 
 data6 <= my_rom(7509); 
 data7 <= my_rom(8864); 
 data8 <= my_rom(10219); 
 data9 <= my_rom(11574); 
 data10 <= my_rom(12929);
when "01011011111" => 
 data1 <= my_rom(735); 
 data2 <= my_rom(2090); 
 data3 <= my_rom(3445); 
 data4 <= my_rom(4800); 
 data5 <= my_rom(6155); 
 data6 <= my_rom(7510); 
 data7 <= my_rom(8865); 
 data8 <= my_rom(10220); 
 data9 <= my_rom(11575); 
 data10 <= my_rom(12930);
when "01011100000" => 
 data1 <= my_rom(736); 
 data2 <= my_rom(2091); 
 data3 <= my_rom(3446); 
 data4 <= my_rom(4801); 
 data5 <= my_rom(6156); 
 data6 <= my_rom(7511); 
 data7 <= my_rom(8866); 
 data8 <= my_rom(10221); 
 data9 <= my_rom(11576); 
 data10 <= my_rom(12931);
when "01011100001" => 
 data1 <= my_rom(737); 
 data2 <= my_rom(2092); 
 data3 <= my_rom(3447); 
 data4 <= my_rom(4802); 
 data5 <= my_rom(6157); 
 data6 <= my_rom(7512); 
 data7 <= my_rom(8867); 
 data8 <= my_rom(10222); 
 data9 <= my_rom(11577); 
 data10 <= my_rom(12932);
when "01011100010" => 
 data1 <= my_rom(738); 
 data2 <= my_rom(2093); 
 data3 <= my_rom(3448); 
 data4 <= my_rom(4803); 
 data5 <= my_rom(6158); 
 data6 <= my_rom(7513); 
 data7 <= my_rom(8868); 
 data8 <= my_rom(10223); 
 data9 <= my_rom(11578); 
 data10 <= my_rom(12933);
when "01011100011" => 
 data1 <= my_rom(739); 
 data2 <= my_rom(2094); 
 data3 <= my_rom(3449); 
 data4 <= my_rom(4804); 
 data5 <= my_rom(6159); 
 data6 <= my_rom(7514); 
 data7 <= my_rom(8869); 
 data8 <= my_rom(10224); 
 data9 <= my_rom(11579); 
 data10 <= my_rom(12934);
when "01011100100" => 
 data1 <= my_rom(740); 
 data2 <= my_rom(2095); 
 data3 <= my_rom(3450); 
 data4 <= my_rom(4805); 
 data5 <= my_rom(6160); 
 data6 <= my_rom(7515); 
 data7 <= my_rom(8870); 
 data8 <= my_rom(10225); 
 data9 <= my_rom(11580); 
 data10 <= my_rom(12935);
when "01011100101" => 
 data1 <= my_rom(741); 
 data2 <= my_rom(2096); 
 data3 <= my_rom(3451); 
 data4 <= my_rom(4806); 
 data5 <= my_rom(6161); 
 data6 <= my_rom(7516); 
 data7 <= my_rom(8871); 
 data8 <= my_rom(10226); 
 data9 <= my_rom(11581); 
 data10 <= my_rom(12936);
when "01011100110" => 
 data1 <= my_rom(742); 
 data2 <= my_rom(2097); 
 data3 <= my_rom(3452); 
 data4 <= my_rom(4807); 
 data5 <= my_rom(6162); 
 data6 <= my_rom(7517); 
 data7 <= my_rom(8872); 
 data8 <= my_rom(10227); 
 data9 <= my_rom(11582); 
 data10 <= my_rom(12937);
when "01011100111" => 
 data1 <= my_rom(743); 
 data2 <= my_rom(2098); 
 data3 <= my_rom(3453); 
 data4 <= my_rom(4808); 
 data5 <= my_rom(6163); 
 data6 <= my_rom(7518); 
 data7 <= my_rom(8873); 
 data8 <= my_rom(10228); 
 data9 <= my_rom(11583); 
 data10 <= my_rom(12938);
when "01011101000" => 
 data1 <= my_rom(744); 
 data2 <= my_rom(2099); 
 data3 <= my_rom(3454); 
 data4 <= my_rom(4809); 
 data5 <= my_rom(6164); 
 data6 <= my_rom(7519); 
 data7 <= my_rom(8874); 
 data8 <= my_rom(10229); 
 data9 <= my_rom(11584); 
 data10 <= my_rom(12939);
when "01011101001" => 
 data1 <= my_rom(745); 
 data2 <= my_rom(2100); 
 data3 <= my_rom(3455); 
 data4 <= my_rom(4810); 
 data5 <= my_rom(6165); 
 data6 <= my_rom(7520); 
 data7 <= my_rom(8875); 
 data8 <= my_rom(10230); 
 data9 <= my_rom(11585); 
 data10 <= my_rom(12940);
when "01011101010" => 
 data1 <= my_rom(746); 
 data2 <= my_rom(2101); 
 data3 <= my_rom(3456); 
 data4 <= my_rom(4811); 
 data5 <= my_rom(6166); 
 data6 <= my_rom(7521); 
 data7 <= my_rom(8876); 
 data8 <= my_rom(10231); 
 data9 <= my_rom(11586); 
 data10 <= my_rom(12941);
when "01011101011" => 
 data1 <= my_rom(747); 
 data2 <= my_rom(2102); 
 data3 <= my_rom(3457); 
 data4 <= my_rom(4812); 
 data5 <= my_rom(6167); 
 data6 <= my_rom(7522); 
 data7 <= my_rom(8877); 
 data8 <= my_rom(10232); 
 data9 <= my_rom(11587); 
 data10 <= my_rom(12942);
when "01011101100" => 
 data1 <= my_rom(748); 
 data2 <= my_rom(2103); 
 data3 <= my_rom(3458); 
 data4 <= my_rom(4813); 
 data5 <= my_rom(6168); 
 data6 <= my_rom(7523); 
 data7 <= my_rom(8878); 
 data8 <= my_rom(10233); 
 data9 <= my_rom(11588); 
 data10 <= my_rom(12943);
when "01011101101" => 
 data1 <= my_rom(749); 
 data2 <= my_rom(2104); 
 data3 <= my_rom(3459); 
 data4 <= my_rom(4814); 
 data5 <= my_rom(6169); 
 data6 <= my_rom(7524); 
 data7 <= my_rom(8879); 
 data8 <= my_rom(10234); 
 data9 <= my_rom(11589); 
 data10 <= my_rom(12944);
when "01011101110" => 
 data1 <= my_rom(750); 
 data2 <= my_rom(2105); 
 data3 <= my_rom(3460); 
 data4 <= my_rom(4815); 
 data5 <= my_rom(6170); 
 data6 <= my_rom(7525); 
 data7 <= my_rom(8880); 
 data8 <= my_rom(10235); 
 data9 <= my_rom(11590); 
 data10 <= my_rom(12945);
when "01011101111" => 
 data1 <= my_rom(751); 
 data2 <= my_rom(2106); 
 data3 <= my_rom(3461); 
 data4 <= my_rom(4816); 
 data5 <= my_rom(6171); 
 data6 <= my_rom(7526); 
 data7 <= my_rom(8881); 
 data8 <= my_rom(10236); 
 data9 <= my_rom(11591); 
 data10 <= my_rom(12946);
when "01011110000" => 
 data1 <= my_rom(752); 
 data2 <= my_rom(2107); 
 data3 <= my_rom(3462); 
 data4 <= my_rom(4817); 
 data5 <= my_rom(6172); 
 data6 <= my_rom(7527); 
 data7 <= my_rom(8882); 
 data8 <= my_rom(10237); 
 data9 <= my_rom(11592); 
 data10 <= my_rom(12947);
when "01011110001" => 
 data1 <= my_rom(753); 
 data2 <= my_rom(2108); 
 data3 <= my_rom(3463); 
 data4 <= my_rom(4818); 
 data5 <= my_rom(6173); 
 data6 <= my_rom(7528); 
 data7 <= my_rom(8883); 
 data8 <= my_rom(10238); 
 data9 <= my_rom(11593); 
 data10 <= my_rom(12948);
when "01011110010" => 
 data1 <= my_rom(754); 
 data2 <= my_rom(2109); 
 data3 <= my_rom(3464); 
 data4 <= my_rom(4819); 
 data5 <= my_rom(6174); 
 data6 <= my_rom(7529); 
 data7 <= my_rom(8884); 
 data8 <= my_rom(10239); 
 data9 <= my_rom(11594); 
 data10 <= my_rom(12949);
when "01011110011" => 
 data1 <= my_rom(755); 
 data2 <= my_rom(2110); 
 data3 <= my_rom(3465); 
 data4 <= my_rom(4820); 
 data5 <= my_rom(6175); 
 data6 <= my_rom(7530); 
 data7 <= my_rom(8885); 
 data8 <= my_rom(10240); 
 data9 <= my_rom(11595); 
 data10 <= my_rom(12950);
when "01011110100" => 
 data1 <= my_rom(756); 
 data2 <= my_rom(2111); 
 data3 <= my_rom(3466); 
 data4 <= my_rom(4821); 
 data5 <= my_rom(6176); 
 data6 <= my_rom(7531); 
 data7 <= my_rom(8886); 
 data8 <= my_rom(10241); 
 data9 <= my_rom(11596); 
 data10 <= my_rom(12951);
when "01011110101" => 
 data1 <= my_rom(757); 
 data2 <= my_rom(2112); 
 data3 <= my_rom(3467); 
 data4 <= my_rom(4822); 
 data5 <= my_rom(6177); 
 data6 <= my_rom(7532); 
 data7 <= my_rom(8887); 
 data8 <= my_rom(10242); 
 data9 <= my_rom(11597); 
 data10 <= my_rom(12952);
when "01011110110" => 
 data1 <= my_rom(758); 
 data2 <= my_rom(2113); 
 data3 <= my_rom(3468); 
 data4 <= my_rom(4823); 
 data5 <= my_rom(6178); 
 data6 <= my_rom(7533); 
 data7 <= my_rom(8888); 
 data8 <= my_rom(10243); 
 data9 <= my_rom(11598); 
 data10 <= my_rom(12953);
when "01011110111" => 
 data1 <= my_rom(759); 
 data2 <= my_rom(2114); 
 data3 <= my_rom(3469); 
 data4 <= my_rom(4824); 
 data5 <= my_rom(6179); 
 data6 <= my_rom(7534); 
 data7 <= my_rom(8889); 
 data8 <= my_rom(10244); 
 data9 <= my_rom(11599); 
 data10 <= my_rom(12954);
when "01011111000" => 
 data1 <= my_rom(760); 
 data2 <= my_rom(2115); 
 data3 <= my_rom(3470); 
 data4 <= my_rom(4825); 
 data5 <= my_rom(6180); 
 data6 <= my_rom(7535); 
 data7 <= my_rom(8890); 
 data8 <= my_rom(10245); 
 data9 <= my_rom(11600); 
 data10 <= my_rom(12955);
when "01011111001" => 
 data1 <= my_rom(761); 
 data2 <= my_rom(2116); 
 data3 <= my_rom(3471); 
 data4 <= my_rom(4826); 
 data5 <= my_rom(6181); 
 data6 <= my_rom(7536); 
 data7 <= my_rom(8891); 
 data8 <= my_rom(10246); 
 data9 <= my_rom(11601); 
 data10 <= my_rom(12956);
when "01011111010" => 
 data1 <= my_rom(762); 
 data2 <= my_rom(2117); 
 data3 <= my_rom(3472); 
 data4 <= my_rom(4827); 
 data5 <= my_rom(6182); 
 data6 <= my_rom(7537); 
 data7 <= my_rom(8892); 
 data8 <= my_rom(10247); 
 data9 <= my_rom(11602); 
 data10 <= my_rom(12957);
when "01011111011" => 
 data1 <= my_rom(763); 
 data2 <= my_rom(2118); 
 data3 <= my_rom(3473); 
 data4 <= my_rom(4828); 
 data5 <= my_rom(6183); 
 data6 <= my_rom(7538); 
 data7 <= my_rom(8893); 
 data8 <= my_rom(10248); 
 data9 <= my_rom(11603); 
 data10 <= my_rom(12958);
when "01011111100" => 
 data1 <= my_rom(764); 
 data2 <= my_rom(2119); 
 data3 <= my_rom(3474); 
 data4 <= my_rom(4829); 
 data5 <= my_rom(6184); 
 data6 <= my_rom(7539); 
 data7 <= my_rom(8894); 
 data8 <= my_rom(10249); 
 data9 <= my_rom(11604); 
 data10 <= my_rom(12959);
when "01011111101" => 
 data1 <= my_rom(765); 
 data2 <= my_rom(2120); 
 data3 <= my_rom(3475); 
 data4 <= my_rom(4830); 
 data5 <= my_rom(6185); 
 data6 <= my_rom(7540); 
 data7 <= my_rom(8895); 
 data8 <= my_rom(10250); 
 data9 <= my_rom(11605); 
 data10 <= my_rom(12960);
when "01011111110" => 
 data1 <= my_rom(766); 
 data2 <= my_rom(2121); 
 data3 <= my_rom(3476); 
 data4 <= my_rom(4831); 
 data5 <= my_rom(6186); 
 data6 <= my_rom(7541); 
 data7 <= my_rom(8896); 
 data8 <= my_rom(10251); 
 data9 <= my_rom(11606); 
 data10 <= my_rom(12961);
when "01011111111" => 
 data1 <= my_rom(767); 
 data2 <= my_rom(2122); 
 data3 <= my_rom(3477); 
 data4 <= my_rom(4832); 
 data5 <= my_rom(6187); 
 data6 <= my_rom(7542); 
 data7 <= my_rom(8897); 
 data8 <= my_rom(10252); 
 data9 <= my_rom(11607); 
 data10 <= my_rom(12962);
when "01100000000" => 
 data1 <= my_rom(768); 
 data2 <= my_rom(2123); 
 data3 <= my_rom(3478); 
 data4 <= my_rom(4833); 
 data5 <= my_rom(6188); 
 data6 <= my_rom(7543); 
 data7 <= my_rom(8898); 
 data8 <= my_rom(10253); 
 data9 <= my_rom(11608); 
 data10 <= my_rom(12963);
when "01100000001" => 
 data1 <= my_rom(769); 
 data2 <= my_rom(2124); 
 data3 <= my_rom(3479); 
 data4 <= my_rom(4834); 
 data5 <= my_rom(6189); 
 data6 <= my_rom(7544); 
 data7 <= my_rom(8899); 
 data8 <= my_rom(10254); 
 data9 <= my_rom(11609); 
 data10 <= my_rom(12964);
when "01100000010" => 
 data1 <= my_rom(770); 
 data2 <= my_rom(2125); 
 data3 <= my_rom(3480); 
 data4 <= my_rom(4835); 
 data5 <= my_rom(6190); 
 data6 <= my_rom(7545); 
 data7 <= my_rom(8900); 
 data8 <= my_rom(10255); 
 data9 <= my_rom(11610); 
 data10 <= my_rom(12965);
when "01100000011" => 
 data1 <= my_rom(771); 
 data2 <= my_rom(2126); 
 data3 <= my_rom(3481); 
 data4 <= my_rom(4836); 
 data5 <= my_rom(6191); 
 data6 <= my_rom(7546); 
 data7 <= my_rom(8901); 
 data8 <= my_rom(10256); 
 data9 <= my_rom(11611); 
 data10 <= my_rom(12966);
when "01100000100" => 
 data1 <= my_rom(772); 
 data2 <= my_rom(2127); 
 data3 <= my_rom(3482); 
 data4 <= my_rom(4837); 
 data5 <= my_rom(6192); 
 data6 <= my_rom(7547); 
 data7 <= my_rom(8902); 
 data8 <= my_rom(10257); 
 data9 <= my_rom(11612); 
 data10 <= my_rom(12967);
when "01100000101" => 
 data1 <= my_rom(773); 
 data2 <= my_rom(2128); 
 data3 <= my_rom(3483); 
 data4 <= my_rom(4838); 
 data5 <= my_rom(6193); 
 data6 <= my_rom(7548); 
 data7 <= my_rom(8903); 
 data8 <= my_rom(10258); 
 data9 <= my_rom(11613); 
 data10 <= my_rom(12968);
when "01100000110" => 
 data1 <= my_rom(774); 
 data2 <= my_rom(2129); 
 data3 <= my_rom(3484); 
 data4 <= my_rom(4839); 
 data5 <= my_rom(6194); 
 data6 <= my_rom(7549); 
 data7 <= my_rom(8904); 
 data8 <= my_rom(10259); 
 data9 <= my_rom(11614); 
 data10 <= my_rom(12969);
when "01100000111" => 
 data1 <= my_rom(775); 
 data2 <= my_rom(2130); 
 data3 <= my_rom(3485); 
 data4 <= my_rom(4840); 
 data5 <= my_rom(6195); 
 data6 <= my_rom(7550); 
 data7 <= my_rom(8905); 
 data8 <= my_rom(10260); 
 data9 <= my_rom(11615); 
 data10 <= my_rom(12970);
when "01100001000" => 
 data1 <= my_rom(776); 
 data2 <= my_rom(2131); 
 data3 <= my_rom(3486); 
 data4 <= my_rom(4841); 
 data5 <= my_rom(6196); 
 data6 <= my_rom(7551); 
 data7 <= my_rom(8906); 
 data8 <= my_rom(10261); 
 data9 <= my_rom(11616); 
 data10 <= my_rom(12971);
when "01100001001" => 
 data1 <= my_rom(777); 
 data2 <= my_rom(2132); 
 data3 <= my_rom(3487); 
 data4 <= my_rom(4842); 
 data5 <= my_rom(6197); 
 data6 <= my_rom(7552); 
 data7 <= my_rom(8907); 
 data8 <= my_rom(10262); 
 data9 <= my_rom(11617); 
 data10 <= my_rom(12972);
when "01100001010" => 
 data1 <= my_rom(778); 
 data2 <= my_rom(2133); 
 data3 <= my_rom(3488); 
 data4 <= my_rom(4843); 
 data5 <= my_rom(6198); 
 data6 <= my_rom(7553); 
 data7 <= my_rom(8908); 
 data8 <= my_rom(10263); 
 data9 <= my_rom(11618); 
 data10 <= my_rom(12973);
when "01100001011" => 
 data1 <= my_rom(779); 
 data2 <= my_rom(2134); 
 data3 <= my_rom(3489); 
 data4 <= my_rom(4844); 
 data5 <= my_rom(6199); 
 data6 <= my_rom(7554); 
 data7 <= my_rom(8909); 
 data8 <= my_rom(10264); 
 data9 <= my_rom(11619); 
 data10 <= my_rom(12974);
when "01100001100" => 
 data1 <= my_rom(780); 
 data2 <= my_rom(2135); 
 data3 <= my_rom(3490); 
 data4 <= my_rom(4845); 
 data5 <= my_rom(6200); 
 data6 <= my_rom(7555); 
 data7 <= my_rom(8910); 
 data8 <= my_rom(10265); 
 data9 <= my_rom(11620); 
 data10 <= my_rom(12975);
when "01100001101" => 
 data1 <= my_rom(781); 
 data2 <= my_rom(2136); 
 data3 <= my_rom(3491); 
 data4 <= my_rom(4846); 
 data5 <= my_rom(6201); 
 data6 <= my_rom(7556); 
 data7 <= my_rom(8911); 
 data8 <= my_rom(10266); 
 data9 <= my_rom(11621); 
 data10 <= my_rom(12976);
when "01100001110" => 
 data1 <= my_rom(782); 
 data2 <= my_rom(2137); 
 data3 <= my_rom(3492); 
 data4 <= my_rom(4847); 
 data5 <= my_rom(6202); 
 data6 <= my_rom(7557); 
 data7 <= my_rom(8912); 
 data8 <= my_rom(10267); 
 data9 <= my_rom(11622); 
 data10 <= my_rom(12977);
when "01100001111" => 
 data1 <= my_rom(783); 
 data2 <= my_rom(2138); 
 data3 <= my_rom(3493); 
 data4 <= my_rom(4848); 
 data5 <= my_rom(6203); 
 data6 <= my_rom(7558); 
 data7 <= my_rom(8913); 
 data8 <= my_rom(10268); 
 data9 <= my_rom(11623); 
 data10 <= my_rom(12978);
when "01100010000" => 
 data1 <= my_rom(784); 
 data2 <= my_rom(2139); 
 data3 <= my_rom(3494); 
 data4 <= my_rom(4849); 
 data5 <= my_rom(6204); 
 data6 <= my_rom(7559); 
 data7 <= my_rom(8914); 
 data8 <= my_rom(10269); 
 data9 <= my_rom(11624); 
 data10 <= my_rom(12979);
when "01100010001" => 
 data1 <= my_rom(785); 
 data2 <= my_rom(2140); 
 data3 <= my_rom(3495); 
 data4 <= my_rom(4850); 
 data5 <= my_rom(6205); 
 data6 <= my_rom(7560); 
 data7 <= my_rom(8915); 
 data8 <= my_rom(10270); 
 data9 <= my_rom(11625); 
 data10 <= my_rom(12980);
when "01100010010" => 
 data1 <= my_rom(786); 
 data2 <= my_rom(2141); 
 data3 <= my_rom(3496); 
 data4 <= my_rom(4851); 
 data5 <= my_rom(6206); 
 data6 <= my_rom(7561); 
 data7 <= my_rom(8916); 
 data8 <= my_rom(10271); 
 data9 <= my_rom(11626); 
 data10 <= my_rom(12981);
when "01100010011" => 
 data1 <= my_rom(787); 
 data2 <= my_rom(2142); 
 data3 <= my_rom(3497); 
 data4 <= my_rom(4852); 
 data5 <= my_rom(6207); 
 data6 <= my_rom(7562); 
 data7 <= my_rom(8917); 
 data8 <= my_rom(10272); 
 data9 <= my_rom(11627); 
 data10 <= my_rom(12982);
when "01100010100" => 
 data1 <= my_rom(788); 
 data2 <= my_rom(2143); 
 data3 <= my_rom(3498); 
 data4 <= my_rom(4853); 
 data5 <= my_rom(6208); 
 data6 <= my_rom(7563); 
 data7 <= my_rom(8918); 
 data8 <= my_rom(10273); 
 data9 <= my_rom(11628); 
 data10 <= my_rom(12983);
when "01100010101" => 
 data1 <= my_rom(789); 
 data2 <= my_rom(2144); 
 data3 <= my_rom(3499); 
 data4 <= my_rom(4854); 
 data5 <= my_rom(6209); 
 data6 <= my_rom(7564); 
 data7 <= my_rom(8919); 
 data8 <= my_rom(10274); 
 data9 <= my_rom(11629); 
 data10 <= my_rom(12984);
when "01100010110" => 
 data1 <= my_rom(790); 
 data2 <= my_rom(2145); 
 data3 <= my_rom(3500); 
 data4 <= my_rom(4855); 
 data5 <= my_rom(6210); 
 data6 <= my_rom(7565); 
 data7 <= my_rom(8920); 
 data8 <= my_rom(10275); 
 data9 <= my_rom(11630); 
 data10 <= my_rom(12985);
when "01100010111" => 
 data1 <= my_rom(791); 
 data2 <= my_rom(2146); 
 data3 <= my_rom(3501); 
 data4 <= my_rom(4856); 
 data5 <= my_rom(6211); 
 data6 <= my_rom(7566); 
 data7 <= my_rom(8921); 
 data8 <= my_rom(10276); 
 data9 <= my_rom(11631); 
 data10 <= my_rom(12986);
when "01100011000" => 
 data1 <= my_rom(792); 
 data2 <= my_rom(2147); 
 data3 <= my_rom(3502); 
 data4 <= my_rom(4857); 
 data5 <= my_rom(6212); 
 data6 <= my_rom(7567); 
 data7 <= my_rom(8922); 
 data8 <= my_rom(10277); 
 data9 <= my_rom(11632); 
 data10 <= my_rom(12987);
when "01100011001" => 
 data1 <= my_rom(793); 
 data2 <= my_rom(2148); 
 data3 <= my_rom(3503); 
 data4 <= my_rom(4858); 
 data5 <= my_rom(6213); 
 data6 <= my_rom(7568); 
 data7 <= my_rom(8923); 
 data8 <= my_rom(10278); 
 data9 <= my_rom(11633); 
 data10 <= my_rom(12988);
when "01100011010" => 
 data1 <= my_rom(794); 
 data2 <= my_rom(2149); 
 data3 <= my_rom(3504); 
 data4 <= my_rom(4859); 
 data5 <= my_rom(6214); 
 data6 <= my_rom(7569); 
 data7 <= my_rom(8924); 
 data8 <= my_rom(10279); 
 data9 <= my_rom(11634); 
 data10 <= my_rom(12989);
when "01100011011" => 
 data1 <= my_rom(795); 
 data2 <= my_rom(2150); 
 data3 <= my_rom(3505); 
 data4 <= my_rom(4860); 
 data5 <= my_rom(6215); 
 data6 <= my_rom(7570); 
 data7 <= my_rom(8925); 
 data8 <= my_rom(10280); 
 data9 <= my_rom(11635); 
 data10 <= my_rom(12990);
when "01100011100" => 
 data1 <= my_rom(796); 
 data2 <= my_rom(2151); 
 data3 <= my_rom(3506); 
 data4 <= my_rom(4861); 
 data5 <= my_rom(6216); 
 data6 <= my_rom(7571); 
 data7 <= my_rom(8926); 
 data8 <= my_rom(10281); 
 data9 <= my_rom(11636); 
 data10 <= my_rom(12991);
when "01100011101" => 
 data1 <= my_rom(797); 
 data2 <= my_rom(2152); 
 data3 <= my_rom(3507); 
 data4 <= my_rom(4862); 
 data5 <= my_rom(6217); 
 data6 <= my_rom(7572); 
 data7 <= my_rom(8927); 
 data8 <= my_rom(10282); 
 data9 <= my_rom(11637); 
 data10 <= my_rom(12992);
when "01100011110" => 
 data1 <= my_rom(798); 
 data2 <= my_rom(2153); 
 data3 <= my_rom(3508); 
 data4 <= my_rom(4863); 
 data5 <= my_rom(6218); 
 data6 <= my_rom(7573); 
 data7 <= my_rom(8928); 
 data8 <= my_rom(10283); 
 data9 <= my_rom(11638); 
 data10 <= my_rom(12993);
when "01100011111" => 
 data1 <= my_rom(799); 
 data2 <= my_rom(2154); 
 data3 <= my_rom(3509); 
 data4 <= my_rom(4864); 
 data5 <= my_rom(6219); 
 data6 <= my_rom(7574); 
 data7 <= my_rom(8929); 
 data8 <= my_rom(10284); 
 data9 <= my_rom(11639); 
 data10 <= my_rom(12994);
when "01100100000" => 
 data1 <= my_rom(800); 
 data2 <= my_rom(2155); 
 data3 <= my_rom(3510); 
 data4 <= my_rom(4865); 
 data5 <= my_rom(6220); 
 data6 <= my_rom(7575); 
 data7 <= my_rom(8930); 
 data8 <= my_rom(10285); 
 data9 <= my_rom(11640); 
 data10 <= my_rom(12995);
when "01100100001" => 
 data1 <= my_rom(801); 
 data2 <= my_rom(2156); 
 data3 <= my_rom(3511); 
 data4 <= my_rom(4866); 
 data5 <= my_rom(6221); 
 data6 <= my_rom(7576); 
 data7 <= my_rom(8931); 
 data8 <= my_rom(10286); 
 data9 <= my_rom(11641); 
 data10 <= my_rom(12996);
when "01100100010" => 
 data1 <= my_rom(802); 
 data2 <= my_rom(2157); 
 data3 <= my_rom(3512); 
 data4 <= my_rom(4867); 
 data5 <= my_rom(6222); 
 data6 <= my_rom(7577); 
 data7 <= my_rom(8932); 
 data8 <= my_rom(10287); 
 data9 <= my_rom(11642); 
 data10 <= my_rom(12997);
when "01100100011" => 
 data1 <= my_rom(803); 
 data2 <= my_rom(2158); 
 data3 <= my_rom(3513); 
 data4 <= my_rom(4868); 
 data5 <= my_rom(6223); 
 data6 <= my_rom(7578); 
 data7 <= my_rom(8933); 
 data8 <= my_rom(10288); 
 data9 <= my_rom(11643); 
 data10 <= my_rom(12998);
when "01100100100" => 
 data1 <= my_rom(804); 
 data2 <= my_rom(2159); 
 data3 <= my_rom(3514); 
 data4 <= my_rom(4869); 
 data5 <= my_rom(6224); 
 data6 <= my_rom(7579); 
 data7 <= my_rom(8934); 
 data8 <= my_rom(10289); 
 data9 <= my_rom(11644); 
 data10 <= my_rom(12999);
when "01100100101" => 
 data1 <= my_rom(805); 
 data2 <= my_rom(2160); 
 data3 <= my_rom(3515); 
 data4 <= my_rom(4870); 
 data5 <= my_rom(6225); 
 data6 <= my_rom(7580); 
 data7 <= my_rom(8935); 
 data8 <= my_rom(10290); 
 data9 <= my_rom(11645); 
 data10 <= my_rom(13000);
when "01100100110" => 
 data1 <= my_rom(806); 
 data2 <= my_rom(2161); 
 data3 <= my_rom(3516); 
 data4 <= my_rom(4871); 
 data5 <= my_rom(6226); 
 data6 <= my_rom(7581); 
 data7 <= my_rom(8936); 
 data8 <= my_rom(10291); 
 data9 <= my_rom(11646); 
 data10 <= my_rom(13001);
when "01100100111" => 
 data1 <= my_rom(807); 
 data2 <= my_rom(2162); 
 data3 <= my_rom(3517); 
 data4 <= my_rom(4872); 
 data5 <= my_rom(6227); 
 data6 <= my_rom(7582); 
 data7 <= my_rom(8937); 
 data8 <= my_rom(10292); 
 data9 <= my_rom(11647); 
 data10 <= my_rom(13002);
when "01100101000" => 
 data1 <= my_rom(808); 
 data2 <= my_rom(2163); 
 data3 <= my_rom(3518); 
 data4 <= my_rom(4873); 
 data5 <= my_rom(6228); 
 data6 <= my_rom(7583); 
 data7 <= my_rom(8938); 
 data8 <= my_rom(10293); 
 data9 <= my_rom(11648); 
 data10 <= my_rom(13003);
when "01100101001" => 
 data1 <= my_rom(809); 
 data2 <= my_rom(2164); 
 data3 <= my_rom(3519); 
 data4 <= my_rom(4874); 
 data5 <= my_rom(6229); 
 data6 <= my_rom(7584); 
 data7 <= my_rom(8939); 
 data8 <= my_rom(10294); 
 data9 <= my_rom(11649); 
 data10 <= my_rom(13004);
when "01100101010" => 
 data1 <= my_rom(810); 
 data2 <= my_rom(2165); 
 data3 <= my_rom(3520); 
 data4 <= my_rom(4875); 
 data5 <= my_rom(6230); 
 data6 <= my_rom(7585); 
 data7 <= my_rom(8940); 
 data8 <= my_rom(10295); 
 data9 <= my_rom(11650); 
 data10 <= my_rom(13005);
when "01100101011" => 
 data1 <= my_rom(811); 
 data2 <= my_rom(2166); 
 data3 <= my_rom(3521); 
 data4 <= my_rom(4876); 
 data5 <= my_rom(6231); 
 data6 <= my_rom(7586); 
 data7 <= my_rom(8941); 
 data8 <= my_rom(10296); 
 data9 <= my_rom(11651); 
 data10 <= my_rom(13006);
when "01100101100" => 
 data1 <= my_rom(812); 
 data2 <= my_rom(2167); 
 data3 <= my_rom(3522); 
 data4 <= my_rom(4877); 
 data5 <= my_rom(6232); 
 data6 <= my_rom(7587); 
 data7 <= my_rom(8942); 
 data8 <= my_rom(10297); 
 data9 <= my_rom(11652); 
 data10 <= my_rom(13007);
when "01100101101" => 
 data1 <= my_rom(813); 
 data2 <= my_rom(2168); 
 data3 <= my_rom(3523); 
 data4 <= my_rom(4878); 
 data5 <= my_rom(6233); 
 data6 <= my_rom(7588); 
 data7 <= my_rom(8943); 
 data8 <= my_rom(10298); 
 data9 <= my_rom(11653); 
 data10 <= my_rom(13008);
when "01100101110" => 
 data1 <= my_rom(814); 
 data2 <= my_rom(2169); 
 data3 <= my_rom(3524); 
 data4 <= my_rom(4879); 
 data5 <= my_rom(6234); 
 data6 <= my_rom(7589); 
 data7 <= my_rom(8944); 
 data8 <= my_rom(10299); 
 data9 <= my_rom(11654); 
 data10 <= my_rom(13009);
when "01100101111" => 
 data1 <= my_rom(815); 
 data2 <= my_rom(2170); 
 data3 <= my_rom(3525); 
 data4 <= my_rom(4880); 
 data5 <= my_rom(6235); 
 data6 <= my_rom(7590); 
 data7 <= my_rom(8945); 
 data8 <= my_rom(10300); 
 data9 <= my_rom(11655); 
 data10 <= my_rom(13010);
when "01100110000" => 
 data1 <= my_rom(816); 
 data2 <= my_rom(2171); 
 data3 <= my_rom(3526); 
 data4 <= my_rom(4881); 
 data5 <= my_rom(6236); 
 data6 <= my_rom(7591); 
 data7 <= my_rom(8946); 
 data8 <= my_rom(10301); 
 data9 <= my_rom(11656); 
 data10 <= my_rom(13011);
when "01100110001" => 
 data1 <= my_rom(817); 
 data2 <= my_rom(2172); 
 data3 <= my_rom(3527); 
 data4 <= my_rom(4882); 
 data5 <= my_rom(6237); 
 data6 <= my_rom(7592); 
 data7 <= my_rom(8947); 
 data8 <= my_rom(10302); 
 data9 <= my_rom(11657); 
 data10 <= my_rom(13012);
when "01100110010" => 
 data1 <= my_rom(818); 
 data2 <= my_rom(2173); 
 data3 <= my_rom(3528); 
 data4 <= my_rom(4883); 
 data5 <= my_rom(6238); 
 data6 <= my_rom(7593); 
 data7 <= my_rom(8948); 
 data8 <= my_rom(10303); 
 data9 <= my_rom(11658); 
 data10 <= my_rom(13013);
when "01100110011" => 
 data1 <= my_rom(819); 
 data2 <= my_rom(2174); 
 data3 <= my_rom(3529); 
 data4 <= my_rom(4884); 
 data5 <= my_rom(6239); 
 data6 <= my_rom(7594); 
 data7 <= my_rom(8949); 
 data8 <= my_rom(10304); 
 data9 <= my_rom(11659); 
 data10 <= my_rom(13014);
when "01100110100" => 
 data1 <= my_rom(820); 
 data2 <= my_rom(2175); 
 data3 <= my_rom(3530); 
 data4 <= my_rom(4885); 
 data5 <= my_rom(6240); 
 data6 <= my_rom(7595); 
 data7 <= my_rom(8950); 
 data8 <= my_rom(10305); 
 data9 <= my_rom(11660); 
 data10 <= my_rom(13015);
when "01100110101" => 
 data1 <= my_rom(821); 
 data2 <= my_rom(2176); 
 data3 <= my_rom(3531); 
 data4 <= my_rom(4886); 
 data5 <= my_rom(6241); 
 data6 <= my_rom(7596); 
 data7 <= my_rom(8951); 
 data8 <= my_rom(10306); 
 data9 <= my_rom(11661); 
 data10 <= my_rom(13016);
when "01100110110" => 
 data1 <= my_rom(822); 
 data2 <= my_rom(2177); 
 data3 <= my_rom(3532); 
 data4 <= my_rom(4887); 
 data5 <= my_rom(6242); 
 data6 <= my_rom(7597); 
 data7 <= my_rom(8952); 
 data8 <= my_rom(10307); 
 data9 <= my_rom(11662); 
 data10 <= my_rom(13017);
when "01100110111" => 
 data1 <= my_rom(823); 
 data2 <= my_rom(2178); 
 data3 <= my_rom(3533); 
 data4 <= my_rom(4888); 
 data5 <= my_rom(6243); 
 data6 <= my_rom(7598); 
 data7 <= my_rom(8953); 
 data8 <= my_rom(10308); 
 data9 <= my_rom(11663); 
 data10 <= my_rom(13018);
when "01100111000" => 
 data1 <= my_rom(824); 
 data2 <= my_rom(2179); 
 data3 <= my_rom(3534); 
 data4 <= my_rom(4889); 
 data5 <= my_rom(6244); 
 data6 <= my_rom(7599); 
 data7 <= my_rom(8954); 
 data8 <= my_rom(10309); 
 data9 <= my_rom(11664); 
 data10 <= my_rom(13019);
when "01100111001" => 
 data1 <= my_rom(825); 
 data2 <= my_rom(2180); 
 data3 <= my_rom(3535); 
 data4 <= my_rom(4890); 
 data5 <= my_rom(6245); 
 data6 <= my_rom(7600); 
 data7 <= my_rom(8955); 
 data8 <= my_rom(10310); 
 data9 <= my_rom(11665); 
 data10 <= my_rom(13020);
when "01100111010" => 
 data1 <= my_rom(826); 
 data2 <= my_rom(2181); 
 data3 <= my_rom(3536); 
 data4 <= my_rom(4891); 
 data5 <= my_rom(6246); 
 data6 <= my_rom(7601); 
 data7 <= my_rom(8956); 
 data8 <= my_rom(10311); 
 data9 <= my_rom(11666); 
 data10 <= my_rom(13021);
when "01100111011" => 
 data1 <= my_rom(827); 
 data2 <= my_rom(2182); 
 data3 <= my_rom(3537); 
 data4 <= my_rom(4892); 
 data5 <= my_rom(6247); 
 data6 <= my_rom(7602); 
 data7 <= my_rom(8957); 
 data8 <= my_rom(10312); 
 data9 <= my_rom(11667); 
 data10 <= my_rom(13022);
when "01100111100" => 
 data1 <= my_rom(828); 
 data2 <= my_rom(2183); 
 data3 <= my_rom(3538); 
 data4 <= my_rom(4893); 
 data5 <= my_rom(6248); 
 data6 <= my_rom(7603); 
 data7 <= my_rom(8958); 
 data8 <= my_rom(10313); 
 data9 <= my_rom(11668); 
 data10 <= my_rom(13023);
when "01100111101" => 
 data1 <= my_rom(829); 
 data2 <= my_rom(2184); 
 data3 <= my_rom(3539); 
 data4 <= my_rom(4894); 
 data5 <= my_rom(6249); 
 data6 <= my_rom(7604); 
 data7 <= my_rom(8959); 
 data8 <= my_rom(10314); 
 data9 <= my_rom(11669); 
 data10 <= my_rom(13024);
when "01100111110" => 
 data1 <= my_rom(830); 
 data2 <= my_rom(2185); 
 data3 <= my_rom(3540); 
 data4 <= my_rom(4895); 
 data5 <= my_rom(6250); 
 data6 <= my_rom(7605); 
 data7 <= my_rom(8960); 
 data8 <= my_rom(10315); 
 data9 <= my_rom(11670); 
 data10 <= my_rom(13025);
when "01100111111" => 
 data1 <= my_rom(831); 
 data2 <= my_rom(2186); 
 data3 <= my_rom(3541); 
 data4 <= my_rom(4896); 
 data5 <= my_rom(6251); 
 data6 <= my_rom(7606); 
 data7 <= my_rom(8961); 
 data8 <= my_rom(10316); 
 data9 <= my_rom(11671); 
 data10 <= my_rom(13026);
when "01101000000" => 
 data1 <= my_rom(832); 
 data2 <= my_rom(2187); 
 data3 <= my_rom(3542); 
 data4 <= my_rom(4897); 
 data5 <= my_rom(6252); 
 data6 <= my_rom(7607); 
 data7 <= my_rom(8962); 
 data8 <= my_rom(10317); 
 data9 <= my_rom(11672); 
 data10 <= my_rom(13027);
when "01101000001" => 
 data1 <= my_rom(833); 
 data2 <= my_rom(2188); 
 data3 <= my_rom(3543); 
 data4 <= my_rom(4898); 
 data5 <= my_rom(6253); 
 data6 <= my_rom(7608); 
 data7 <= my_rom(8963); 
 data8 <= my_rom(10318); 
 data9 <= my_rom(11673); 
 data10 <= my_rom(13028);
when "01101000010" => 
 data1 <= my_rom(834); 
 data2 <= my_rom(2189); 
 data3 <= my_rom(3544); 
 data4 <= my_rom(4899); 
 data5 <= my_rom(6254); 
 data6 <= my_rom(7609); 
 data7 <= my_rom(8964); 
 data8 <= my_rom(10319); 
 data9 <= my_rom(11674); 
 data10 <= my_rom(13029);
when "01101000011" => 
 data1 <= my_rom(835); 
 data2 <= my_rom(2190); 
 data3 <= my_rom(3545); 
 data4 <= my_rom(4900); 
 data5 <= my_rom(6255); 
 data6 <= my_rom(7610); 
 data7 <= my_rom(8965); 
 data8 <= my_rom(10320); 
 data9 <= my_rom(11675); 
 data10 <= my_rom(13030);
when "01101000100" => 
 data1 <= my_rom(836); 
 data2 <= my_rom(2191); 
 data3 <= my_rom(3546); 
 data4 <= my_rom(4901); 
 data5 <= my_rom(6256); 
 data6 <= my_rom(7611); 
 data7 <= my_rom(8966); 
 data8 <= my_rom(10321); 
 data9 <= my_rom(11676); 
 data10 <= my_rom(13031);
when "01101000101" => 
 data1 <= my_rom(837); 
 data2 <= my_rom(2192); 
 data3 <= my_rom(3547); 
 data4 <= my_rom(4902); 
 data5 <= my_rom(6257); 
 data6 <= my_rom(7612); 
 data7 <= my_rom(8967); 
 data8 <= my_rom(10322); 
 data9 <= my_rom(11677); 
 data10 <= my_rom(13032);
when "01101000110" => 
 data1 <= my_rom(838); 
 data2 <= my_rom(2193); 
 data3 <= my_rom(3548); 
 data4 <= my_rom(4903); 
 data5 <= my_rom(6258); 
 data6 <= my_rom(7613); 
 data7 <= my_rom(8968); 
 data8 <= my_rom(10323); 
 data9 <= my_rom(11678); 
 data10 <= my_rom(13033);
when "01101000111" => 
 data1 <= my_rom(839); 
 data2 <= my_rom(2194); 
 data3 <= my_rom(3549); 
 data4 <= my_rom(4904); 
 data5 <= my_rom(6259); 
 data6 <= my_rom(7614); 
 data7 <= my_rom(8969); 
 data8 <= my_rom(10324); 
 data9 <= my_rom(11679); 
 data10 <= my_rom(13034);
when "01101001000" => 
 data1 <= my_rom(840); 
 data2 <= my_rom(2195); 
 data3 <= my_rom(3550); 
 data4 <= my_rom(4905); 
 data5 <= my_rom(6260); 
 data6 <= my_rom(7615); 
 data7 <= my_rom(8970); 
 data8 <= my_rom(10325); 
 data9 <= my_rom(11680); 
 data10 <= my_rom(13035);
when "01101001001" => 
 data1 <= my_rom(841); 
 data2 <= my_rom(2196); 
 data3 <= my_rom(3551); 
 data4 <= my_rom(4906); 
 data5 <= my_rom(6261); 
 data6 <= my_rom(7616); 
 data7 <= my_rom(8971); 
 data8 <= my_rom(10326); 
 data9 <= my_rom(11681); 
 data10 <= my_rom(13036);
when "01101001010" => 
 data1 <= my_rom(842); 
 data2 <= my_rom(2197); 
 data3 <= my_rom(3552); 
 data4 <= my_rom(4907); 
 data5 <= my_rom(6262); 
 data6 <= my_rom(7617); 
 data7 <= my_rom(8972); 
 data8 <= my_rom(10327); 
 data9 <= my_rom(11682); 
 data10 <= my_rom(13037);
when "01101001011" => 
 data1 <= my_rom(843); 
 data2 <= my_rom(2198); 
 data3 <= my_rom(3553); 
 data4 <= my_rom(4908); 
 data5 <= my_rom(6263); 
 data6 <= my_rom(7618); 
 data7 <= my_rom(8973); 
 data8 <= my_rom(10328); 
 data9 <= my_rom(11683); 
 data10 <= my_rom(13038);
when "01101001100" => 
 data1 <= my_rom(844); 
 data2 <= my_rom(2199); 
 data3 <= my_rom(3554); 
 data4 <= my_rom(4909); 
 data5 <= my_rom(6264); 
 data6 <= my_rom(7619); 
 data7 <= my_rom(8974); 
 data8 <= my_rom(10329); 
 data9 <= my_rom(11684); 
 data10 <= my_rom(13039);
when "01101001101" => 
 data1 <= my_rom(845); 
 data2 <= my_rom(2200); 
 data3 <= my_rom(3555); 
 data4 <= my_rom(4910); 
 data5 <= my_rom(6265); 
 data6 <= my_rom(7620); 
 data7 <= my_rom(8975); 
 data8 <= my_rom(10330); 
 data9 <= my_rom(11685); 
 data10 <= my_rom(13040);
when "01101001110" => 
 data1 <= my_rom(846); 
 data2 <= my_rom(2201); 
 data3 <= my_rom(3556); 
 data4 <= my_rom(4911); 
 data5 <= my_rom(6266); 
 data6 <= my_rom(7621); 
 data7 <= my_rom(8976); 
 data8 <= my_rom(10331); 
 data9 <= my_rom(11686); 
 data10 <= my_rom(13041);
when "01101001111" => 
 data1 <= my_rom(847); 
 data2 <= my_rom(2202); 
 data3 <= my_rom(3557); 
 data4 <= my_rom(4912); 
 data5 <= my_rom(6267); 
 data6 <= my_rom(7622); 
 data7 <= my_rom(8977); 
 data8 <= my_rom(10332); 
 data9 <= my_rom(11687); 
 data10 <= my_rom(13042);
when "01101010000" => 
 data1 <= my_rom(848); 
 data2 <= my_rom(2203); 
 data3 <= my_rom(3558); 
 data4 <= my_rom(4913); 
 data5 <= my_rom(6268); 
 data6 <= my_rom(7623); 
 data7 <= my_rom(8978); 
 data8 <= my_rom(10333); 
 data9 <= my_rom(11688); 
 data10 <= my_rom(13043);
when "01101010001" => 
 data1 <= my_rom(849); 
 data2 <= my_rom(2204); 
 data3 <= my_rom(3559); 
 data4 <= my_rom(4914); 
 data5 <= my_rom(6269); 
 data6 <= my_rom(7624); 
 data7 <= my_rom(8979); 
 data8 <= my_rom(10334); 
 data9 <= my_rom(11689); 
 data10 <= my_rom(13044);
when "01101010010" => 
 data1 <= my_rom(850); 
 data2 <= my_rom(2205); 
 data3 <= my_rom(3560); 
 data4 <= my_rom(4915); 
 data5 <= my_rom(6270); 
 data6 <= my_rom(7625); 
 data7 <= my_rom(8980); 
 data8 <= my_rom(10335); 
 data9 <= my_rom(11690); 
 data10 <= my_rom(13045);
when "01101010011" => 
 data1 <= my_rom(851); 
 data2 <= my_rom(2206); 
 data3 <= my_rom(3561); 
 data4 <= my_rom(4916); 
 data5 <= my_rom(6271); 
 data6 <= my_rom(7626); 
 data7 <= my_rom(8981); 
 data8 <= my_rom(10336); 
 data9 <= my_rom(11691); 
 data10 <= my_rom(13046);
when "01101010100" => 
 data1 <= my_rom(852); 
 data2 <= my_rom(2207); 
 data3 <= my_rom(3562); 
 data4 <= my_rom(4917); 
 data5 <= my_rom(6272); 
 data6 <= my_rom(7627); 
 data7 <= my_rom(8982); 
 data8 <= my_rom(10337); 
 data9 <= my_rom(11692); 
 data10 <= my_rom(13047);
when "01101010101" => 
 data1 <= my_rom(853); 
 data2 <= my_rom(2208); 
 data3 <= my_rom(3563); 
 data4 <= my_rom(4918); 
 data5 <= my_rom(6273); 
 data6 <= my_rom(7628); 
 data7 <= my_rom(8983); 
 data8 <= my_rom(10338); 
 data9 <= my_rom(11693); 
 data10 <= my_rom(13048);
when "01101010110" => 
 data1 <= my_rom(854); 
 data2 <= my_rom(2209); 
 data3 <= my_rom(3564); 
 data4 <= my_rom(4919); 
 data5 <= my_rom(6274); 
 data6 <= my_rom(7629); 
 data7 <= my_rom(8984); 
 data8 <= my_rom(10339); 
 data9 <= my_rom(11694); 
 data10 <= my_rom(13049);
when "01101010111" => 
 data1 <= my_rom(855); 
 data2 <= my_rom(2210); 
 data3 <= my_rom(3565); 
 data4 <= my_rom(4920); 
 data5 <= my_rom(6275); 
 data6 <= my_rom(7630); 
 data7 <= my_rom(8985); 
 data8 <= my_rom(10340); 
 data9 <= my_rom(11695); 
 data10 <= my_rom(13050);
when "01101011000" => 
 data1 <= my_rom(856); 
 data2 <= my_rom(2211); 
 data3 <= my_rom(3566); 
 data4 <= my_rom(4921); 
 data5 <= my_rom(6276); 
 data6 <= my_rom(7631); 
 data7 <= my_rom(8986); 
 data8 <= my_rom(10341); 
 data9 <= my_rom(11696); 
 data10 <= my_rom(13051);
when "01101011001" => 
 data1 <= my_rom(857); 
 data2 <= my_rom(2212); 
 data3 <= my_rom(3567); 
 data4 <= my_rom(4922); 
 data5 <= my_rom(6277); 
 data6 <= my_rom(7632); 
 data7 <= my_rom(8987); 
 data8 <= my_rom(10342); 
 data9 <= my_rom(11697); 
 data10 <= my_rom(13052);
when "01101011010" => 
 data1 <= my_rom(858); 
 data2 <= my_rom(2213); 
 data3 <= my_rom(3568); 
 data4 <= my_rom(4923); 
 data5 <= my_rom(6278); 
 data6 <= my_rom(7633); 
 data7 <= my_rom(8988); 
 data8 <= my_rom(10343); 
 data9 <= my_rom(11698); 
 data10 <= my_rom(13053);
when "01101011011" => 
 data1 <= my_rom(859); 
 data2 <= my_rom(2214); 
 data3 <= my_rom(3569); 
 data4 <= my_rom(4924); 
 data5 <= my_rom(6279); 
 data6 <= my_rom(7634); 
 data7 <= my_rom(8989); 
 data8 <= my_rom(10344); 
 data9 <= my_rom(11699); 
 data10 <= my_rom(13054);
when "01101011100" => 
 data1 <= my_rom(860); 
 data2 <= my_rom(2215); 
 data3 <= my_rom(3570); 
 data4 <= my_rom(4925); 
 data5 <= my_rom(6280); 
 data6 <= my_rom(7635); 
 data7 <= my_rom(8990); 
 data8 <= my_rom(10345); 
 data9 <= my_rom(11700); 
 data10 <= my_rom(13055);
when "01101011101" => 
 data1 <= my_rom(861); 
 data2 <= my_rom(2216); 
 data3 <= my_rom(3571); 
 data4 <= my_rom(4926); 
 data5 <= my_rom(6281); 
 data6 <= my_rom(7636); 
 data7 <= my_rom(8991); 
 data8 <= my_rom(10346); 
 data9 <= my_rom(11701); 
 data10 <= my_rom(13056);
when "01101011110" => 
 data1 <= my_rom(862); 
 data2 <= my_rom(2217); 
 data3 <= my_rom(3572); 
 data4 <= my_rom(4927); 
 data5 <= my_rom(6282); 
 data6 <= my_rom(7637); 
 data7 <= my_rom(8992); 
 data8 <= my_rom(10347); 
 data9 <= my_rom(11702); 
 data10 <= my_rom(13057);
when "01101011111" => 
 data1 <= my_rom(863); 
 data2 <= my_rom(2218); 
 data3 <= my_rom(3573); 
 data4 <= my_rom(4928); 
 data5 <= my_rom(6283); 
 data6 <= my_rom(7638); 
 data7 <= my_rom(8993); 
 data8 <= my_rom(10348); 
 data9 <= my_rom(11703); 
 data10 <= my_rom(13058);
when "01101100000" => 
 data1 <= my_rom(864); 
 data2 <= my_rom(2219); 
 data3 <= my_rom(3574); 
 data4 <= my_rom(4929); 
 data5 <= my_rom(6284); 
 data6 <= my_rom(7639); 
 data7 <= my_rom(8994); 
 data8 <= my_rom(10349); 
 data9 <= my_rom(11704); 
 data10 <= my_rom(13059);
when "01101100001" => 
 data1 <= my_rom(865); 
 data2 <= my_rom(2220); 
 data3 <= my_rom(3575); 
 data4 <= my_rom(4930); 
 data5 <= my_rom(6285); 
 data6 <= my_rom(7640); 
 data7 <= my_rom(8995); 
 data8 <= my_rom(10350); 
 data9 <= my_rom(11705); 
 data10 <= my_rom(13060);
when "01101100010" => 
 data1 <= my_rom(866); 
 data2 <= my_rom(2221); 
 data3 <= my_rom(3576); 
 data4 <= my_rom(4931); 
 data5 <= my_rom(6286); 
 data6 <= my_rom(7641); 
 data7 <= my_rom(8996); 
 data8 <= my_rom(10351); 
 data9 <= my_rom(11706); 
 data10 <= my_rom(13061);
when "01101100011" => 
 data1 <= my_rom(867); 
 data2 <= my_rom(2222); 
 data3 <= my_rom(3577); 
 data4 <= my_rom(4932); 
 data5 <= my_rom(6287); 
 data6 <= my_rom(7642); 
 data7 <= my_rom(8997); 
 data8 <= my_rom(10352); 
 data9 <= my_rom(11707); 
 data10 <= my_rom(13062);
when "01101100100" => 
 data1 <= my_rom(868); 
 data2 <= my_rom(2223); 
 data3 <= my_rom(3578); 
 data4 <= my_rom(4933); 
 data5 <= my_rom(6288); 
 data6 <= my_rom(7643); 
 data7 <= my_rom(8998); 
 data8 <= my_rom(10353); 
 data9 <= my_rom(11708); 
 data10 <= my_rom(13063);
when "01101100101" => 
 data1 <= my_rom(869); 
 data2 <= my_rom(2224); 
 data3 <= my_rom(3579); 
 data4 <= my_rom(4934); 
 data5 <= my_rom(6289); 
 data6 <= my_rom(7644); 
 data7 <= my_rom(8999); 
 data8 <= my_rom(10354); 
 data9 <= my_rom(11709); 
 data10 <= my_rom(13064);
when "01101100110" => 
 data1 <= my_rom(870); 
 data2 <= my_rom(2225); 
 data3 <= my_rom(3580); 
 data4 <= my_rom(4935); 
 data5 <= my_rom(6290); 
 data6 <= my_rom(7645); 
 data7 <= my_rom(9000); 
 data8 <= my_rom(10355); 
 data9 <= my_rom(11710); 
 data10 <= my_rom(13065);
when "01101100111" => 
 data1 <= my_rom(871); 
 data2 <= my_rom(2226); 
 data3 <= my_rom(3581); 
 data4 <= my_rom(4936); 
 data5 <= my_rom(6291); 
 data6 <= my_rom(7646); 
 data7 <= my_rom(9001); 
 data8 <= my_rom(10356); 
 data9 <= my_rom(11711); 
 data10 <= my_rom(13066);
when "01101101000" => 
 data1 <= my_rom(872); 
 data2 <= my_rom(2227); 
 data3 <= my_rom(3582); 
 data4 <= my_rom(4937); 
 data5 <= my_rom(6292); 
 data6 <= my_rom(7647); 
 data7 <= my_rom(9002); 
 data8 <= my_rom(10357); 
 data9 <= my_rom(11712); 
 data10 <= my_rom(13067);
when "01101101001" => 
 data1 <= my_rom(873); 
 data2 <= my_rom(2228); 
 data3 <= my_rom(3583); 
 data4 <= my_rom(4938); 
 data5 <= my_rom(6293); 
 data6 <= my_rom(7648); 
 data7 <= my_rom(9003); 
 data8 <= my_rom(10358); 
 data9 <= my_rom(11713); 
 data10 <= my_rom(13068);
when "01101101010" => 
 data1 <= my_rom(874); 
 data2 <= my_rom(2229); 
 data3 <= my_rom(3584); 
 data4 <= my_rom(4939); 
 data5 <= my_rom(6294); 
 data6 <= my_rom(7649); 
 data7 <= my_rom(9004); 
 data8 <= my_rom(10359); 
 data9 <= my_rom(11714); 
 data10 <= my_rom(13069);
when "01101101011" => 
 data1 <= my_rom(875); 
 data2 <= my_rom(2230); 
 data3 <= my_rom(3585); 
 data4 <= my_rom(4940); 
 data5 <= my_rom(6295); 
 data6 <= my_rom(7650); 
 data7 <= my_rom(9005); 
 data8 <= my_rom(10360); 
 data9 <= my_rom(11715); 
 data10 <= my_rom(13070);
when "01101101100" => 
 data1 <= my_rom(876); 
 data2 <= my_rom(2231); 
 data3 <= my_rom(3586); 
 data4 <= my_rom(4941); 
 data5 <= my_rom(6296); 
 data6 <= my_rom(7651); 
 data7 <= my_rom(9006); 
 data8 <= my_rom(10361); 
 data9 <= my_rom(11716); 
 data10 <= my_rom(13071);
when "01101101101" => 
 data1 <= my_rom(877); 
 data2 <= my_rom(2232); 
 data3 <= my_rom(3587); 
 data4 <= my_rom(4942); 
 data5 <= my_rom(6297); 
 data6 <= my_rom(7652); 
 data7 <= my_rom(9007); 
 data8 <= my_rom(10362); 
 data9 <= my_rom(11717); 
 data10 <= my_rom(13072);
when "01101101110" => 
 data1 <= my_rom(878); 
 data2 <= my_rom(2233); 
 data3 <= my_rom(3588); 
 data4 <= my_rom(4943); 
 data5 <= my_rom(6298); 
 data6 <= my_rom(7653); 
 data7 <= my_rom(9008); 
 data8 <= my_rom(10363); 
 data9 <= my_rom(11718); 
 data10 <= my_rom(13073);
when "01101101111" => 
 data1 <= my_rom(879); 
 data2 <= my_rom(2234); 
 data3 <= my_rom(3589); 
 data4 <= my_rom(4944); 
 data5 <= my_rom(6299); 
 data6 <= my_rom(7654); 
 data7 <= my_rom(9009); 
 data8 <= my_rom(10364); 
 data9 <= my_rom(11719); 
 data10 <= my_rom(13074);
when "01101110000" => 
 data1 <= my_rom(880); 
 data2 <= my_rom(2235); 
 data3 <= my_rom(3590); 
 data4 <= my_rom(4945); 
 data5 <= my_rom(6300); 
 data6 <= my_rom(7655); 
 data7 <= my_rom(9010); 
 data8 <= my_rom(10365); 
 data9 <= my_rom(11720); 
 data10 <= my_rom(13075);
when "01101110001" => 
 data1 <= my_rom(881); 
 data2 <= my_rom(2236); 
 data3 <= my_rom(3591); 
 data4 <= my_rom(4946); 
 data5 <= my_rom(6301); 
 data6 <= my_rom(7656); 
 data7 <= my_rom(9011); 
 data8 <= my_rom(10366); 
 data9 <= my_rom(11721); 
 data10 <= my_rom(13076);
when "01101110010" => 
 data1 <= my_rom(882); 
 data2 <= my_rom(2237); 
 data3 <= my_rom(3592); 
 data4 <= my_rom(4947); 
 data5 <= my_rom(6302); 
 data6 <= my_rom(7657); 
 data7 <= my_rom(9012); 
 data8 <= my_rom(10367); 
 data9 <= my_rom(11722); 
 data10 <= my_rom(13077);
when "01101110011" => 
 data1 <= my_rom(883); 
 data2 <= my_rom(2238); 
 data3 <= my_rom(3593); 
 data4 <= my_rom(4948); 
 data5 <= my_rom(6303); 
 data6 <= my_rom(7658); 
 data7 <= my_rom(9013); 
 data8 <= my_rom(10368); 
 data9 <= my_rom(11723); 
 data10 <= my_rom(13078);
when "01101110100" => 
 data1 <= my_rom(884); 
 data2 <= my_rom(2239); 
 data3 <= my_rom(3594); 
 data4 <= my_rom(4949); 
 data5 <= my_rom(6304); 
 data6 <= my_rom(7659); 
 data7 <= my_rom(9014); 
 data8 <= my_rom(10369); 
 data9 <= my_rom(11724); 
 data10 <= my_rom(13079);
when "01101110101" => 
 data1 <= my_rom(885); 
 data2 <= my_rom(2240); 
 data3 <= my_rom(3595); 
 data4 <= my_rom(4950); 
 data5 <= my_rom(6305); 
 data6 <= my_rom(7660); 
 data7 <= my_rom(9015); 
 data8 <= my_rom(10370); 
 data9 <= my_rom(11725); 
 data10 <= my_rom(13080);
when "01101110110" => 
 data1 <= my_rom(886); 
 data2 <= my_rom(2241); 
 data3 <= my_rom(3596); 
 data4 <= my_rom(4951); 
 data5 <= my_rom(6306); 
 data6 <= my_rom(7661); 
 data7 <= my_rom(9016); 
 data8 <= my_rom(10371); 
 data9 <= my_rom(11726); 
 data10 <= my_rom(13081);
when "01101110111" => 
 data1 <= my_rom(887); 
 data2 <= my_rom(2242); 
 data3 <= my_rom(3597); 
 data4 <= my_rom(4952); 
 data5 <= my_rom(6307); 
 data6 <= my_rom(7662); 
 data7 <= my_rom(9017); 
 data8 <= my_rom(10372); 
 data9 <= my_rom(11727); 
 data10 <= my_rom(13082);
when "01101111000" => 
 data1 <= my_rom(888); 
 data2 <= my_rom(2243); 
 data3 <= my_rom(3598); 
 data4 <= my_rom(4953); 
 data5 <= my_rom(6308); 
 data6 <= my_rom(7663); 
 data7 <= my_rom(9018); 
 data8 <= my_rom(10373); 
 data9 <= my_rom(11728); 
 data10 <= my_rom(13083);
when "01101111001" => 
 data1 <= my_rom(889); 
 data2 <= my_rom(2244); 
 data3 <= my_rom(3599); 
 data4 <= my_rom(4954); 
 data5 <= my_rom(6309); 
 data6 <= my_rom(7664); 
 data7 <= my_rom(9019); 
 data8 <= my_rom(10374); 
 data9 <= my_rom(11729); 
 data10 <= my_rom(13084);
when "01101111010" => 
 data1 <= my_rom(890); 
 data2 <= my_rom(2245); 
 data3 <= my_rom(3600); 
 data4 <= my_rom(4955); 
 data5 <= my_rom(6310); 
 data6 <= my_rom(7665); 
 data7 <= my_rom(9020); 
 data8 <= my_rom(10375); 
 data9 <= my_rom(11730); 
 data10 <= my_rom(13085);
when "01101111011" => 
 data1 <= my_rom(891); 
 data2 <= my_rom(2246); 
 data3 <= my_rom(3601); 
 data4 <= my_rom(4956); 
 data5 <= my_rom(6311); 
 data6 <= my_rom(7666); 
 data7 <= my_rom(9021); 
 data8 <= my_rom(10376); 
 data9 <= my_rom(11731); 
 data10 <= my_rom(13086);
when "01101111100" => 
 data1 <= my_rom(892); 
 data2 <= my_rom(2247); 
 data3 <= my_rom(3602); 
 data4 <= my_rom(4957); 
 data5 <= my_rom(6312); 
 data6 <= my_rom(7667); 
 data7 <= my_rom(9022); 
 data8 <= my_rom(10377); 
 data9 <= my_rom(11732); 
 data10 <= my_rom(13087);
when "01101111101" => 
 data1 <= my_rom(893); 
 data2 <= my_rom(2248); 
 data3 <= my_rom(3603); 
 data4 <= my_rom(4958); 
 data5 <= my_rom(6313); 
 data6 <= my_rom(7668); 
 data7 <= my_rom(9023); 
 data8 <= my_rom(10378); 
 data9 <= my_rom(11733); 
 data10 <= my_rom(13088);
when "01101111110" => 
 data1 <= my_rom(894); 
 data2 <= my_rom(2249); 
 data3 <= my_rom(3604); 
 data4 <= my_rom(4959); 
 data5 <= my_rom(6314); 
 data6 <= my_rom(7669); 
 data7 <= my_rom(9024); 
 data8 <= my_rom(10379); 
 data9 <= my_rom(11734); 
 data10 <= my_rom(13089);
when "01101111111" => 
 data1 <= my_rom(895); 
 data2 <= my_rom(2250); 
 data3 <= my_rom(3605); 
 data4 <= my_rom(4960); 
 data5 <= my_rom(6315); 
 data6 <= my_rom(7670); 
 data7 <= my_rom(9025); 
 data8 <= my_rom(10380); 
 data9 <= my_rom(11735); 
 data10 <= my_rom(13090);
when "01110000000" => 
 data1 <= my_rom(896); 
 data2 <= my_rom(2251); 
 data3 <= my_rom(3606); 
 data4 <= my_rom(4961); 
 data5 <= my_rom(6316); 
 data6 <= my_rom(7671); 
 data7 <= my_rom(9026); 
 data8 <= my_rom(10381); 
 data9 <= my_rom(11736); 
 data10 <= my_rom(13091);
when "01110000001" => 
 data1 <= my_rom(897); 
 data2 <= my_rom(2252); 
 data3 <= my_rom(3607); 
 data4 <= my_rom(4962); 
 data5 <= my_rom(6317); 
 data6 <= my_rom(7672); 
 data7 <= my_rom(9027); 
 data8 <= my_rom(10382); 
 data9 <= my_rom(11737); 
 data10 <= my_rom(13092);
when "01110000010" => 
 data1 <= my_rom(898); 
 data2 <= my_rom(2253); 
 data3 <= my_rom(3608); 
 data4 <= my_rom(4963); 
 data5 <= my_rom(6318); 
 data6 <= my_rom(7673); 
 data7 <= my_rom(9028); 
 data8 <= my_rom(10383); 
 data9 <= my_rom(11738); 
 data10 <= my_rom(13093);
when "01110000011" => 
 data1 <= my_rom(899); 
 data2 <= my_rom(2254); 
 data3 <= my_rom(3609); 
 data4 <= my_rom(4964); 
 data5 <= my_rom(6319); 
 data6 <= my_rom(7674); 
 data7 <= my_rom(9029); 
 data8 <= my_rom(10384); 
 data9 <= my_rom(11739); 
 data10 <= my_rom(13094);
when "01110000100" => 
 data1 <= my_rom(900); 
 data2 <= my_rom(2255); 
 data3 <= my_rom(3610); 
 data4 <= my_rom(4965); 
 data5 <= my_rom(6320); 
 data6 <= my_rom(7675); 
 data7 <= my_rom(9030); 
 data8 <= my_rom(10385); 
 data9 <= my_rom(11740); 
 data10 <= my_rom(13095);
when "01110000101" => 
 data1 <= my_rom(901); 
 data2 <= my_rom(2256); 
 data3 <= my_rom(3611); 
 data4 <= my_rom(4966); 
 data5 <= my_rom(6321); 
 data6 <= my_rom(7676); 
 data7 <= my_rom(9031); 
 data8 <= my_rom(10386); 
 data9 <= my_rom(11741); 
 data10 <= my_rom(13096);
when "01110000110" => 
 data1 <= my_rom(902); 
 data2 <= my_rom(2257); 
 data3 <= my_rom(3612); 
 data4 <= my_rom(4967); 
 data5 <= my_rom(6322); 
 data6 <= my_rom(7677); 
 data7 <= my_rom(9032); 
 data8 <= my_rom(10387); 
 data9 <= my_rom(11742); 
 data10 <= my_rom(13097);
when "01110000111" => 
 data1 <= my_rom(903); 
 data2 <= my_rom(2258); 
 data3 <= my_rom(3613); 
 data4 <= my_rom(4968); 
 data5 <= my_rom(6323); 
 data6 <= my_rom(7678); 
 data7 <= my_rom(9033); 
 data8 <= my_rom(10388); 
 data9 <= my_rom(11743); 
 data10 <= my_rom(13098);
when "01110001000" => 
 data1 <= my_rom(904); 
 data2 <= my_rom(2259); 
 data3 <= my_rom(3614); 
 data4 <= my_rom(4969); 
 data5 <= my_rom(6324); 
 data6 <= my_rom(7679); 
 data7 <= my_rom(9034); 
 data8 <= my_rom(10389); 
 data9 <= my_rom(11744); 
 data10 <= my_rom(13099);
when "01110001001" => 
 data1 <= my_rom(905); 
 data2 <= my_rom(2260); 
 data3 <= my_rom(3615); 
 data4 <= my_rom(4970); 
 data5 <= my_rom(6325); 
 data6 <= my_rom(7680); 
 data7 <= my_rom(9035); 
 data8 <= my_rom(10390); 
 data9 <= my_rom(11745); 
 data10 <= my_rom(13100);
when "01110001010" => 
 data1 <= my_rom(906); 
 data2 <= my_rom(2261); 
 data3 <= my_rom(3616); 
 data4 <= my_rom(4971); 
 data5 <= my_rom(6326); 
 data6 <= my_rom(7681); 
 data7 <= my_rom(9036); 
 data8 <= my_rom(10391); 
 data9 <= my_rom(11746); 
 data10 <= my_rom(13101);
when "01110001011" => 
 data1 <= my_rom(907); 
 data2 <= my_rom(2262); 
 data3 <= my_rom(3617); 
 data4 <= my_rom(4972); 
 data5 <= my_rom(6327); 
 data6 <= my_rom(7682); 
 data7 <= my_rom(9037); 
 data8 <= my_rom(10392); 
 data9 <= my_rom(11747); 
 data10 <= my_rom(13102);
when "01110001100" => 
 data1 <= my_rom(908); 
 data2 <= my_rom(2263); 
 data3 <= my_rom(3618); 
 data4 <= my_rom(4973); 
 data5 <= my_rom(6328); 
 data6 <= my_rom(7683); 
 data7 <= my_rom(9038); 
 data8 <= my_rom(10393); 
 data9 <= my_rom(11748); 
 data10 <= my_rom(13103);
when "01110001101" => 
 data1 <= my_rom(909); 
 data2 <= my_rom(2264); 
 data3 <= my_rom(3619); 
 data4 <= my_rom(4974); 
 data5 <= my_rom(6329); 
 data6 <= my_rom(7684); 
 data7 <= my_rom(9039); 
 data8 <= my_rom(10394); 
 data9 <= my_rom(11749); 
 data10 <= my_rom(13104);
when "01110001110" => 
 data1 <= my_rom(910); 
 data2 <= my_rom(2265); 
 data3 <= my_rom(3620); 
 data4 <= my_rom(4975); 
 data5 <= my_rom(6330); 
 data6 <= my_rom(7685); 
 data7 <= my_rom(9040); 
 data8 <= my_rom(10395); 
 data9 <= my_rom(11750); 
 data10 <= my_rom(13105);
when "01110001111" => 
 data1 <= my_rom(911); 
 data2 <= my_rom(2266); 
 data3 <= my_rom(3621); 
 data4 <= my_rom(4976); 
 data5 <= my_rom(6331); 
 data6 <= my_rom(7686); 
 data7 <= my_rom(9041); 
 data8 <= my_rom(10396); 
 data9 <= my_rom(11751); 
 data10 <= my_rom(13106);
when "01110010000" => 
 data1 <= my_rom(912); 
 data2 <= my_rom(2267); 
 data3 <= my_rom(3622); 
 data4 <= my_rom(4977); 
 data5 <= my_rom(6332); 
 data6 <= my_rom(7687); 
 data7 <= my_rom(9042); 
 data8 <= my_rom(10397); 
 data9 <= my_rom(11752); 
 data10 <= my_rom(13107);
when "01110010001" => 
 data1 <= my_rom(913); 
 data2 <= my_rom(2268); 
 data3 <= my_rom(3623); 
 data4 <= my_rom(4978); 
 data5 <= my_rom(6333); 
 data6 <= my_rom(7688); 
 data7 <= my_rom(9043); 
 data8 <= my_rom(10398); 
 data9 <= my_rom(11753); 
 data10 <= my_rom(13108);
when "01110010010" => 
 data1 <= my_rom(914); 
 data2 <= my_rom(2269); 
 data3 <= my_rom(3624); 
 data4 <= my_rom(4979); 
 data5 <= my_rom(6334); 
 data6 <= my_rom(7689); 
 data7 <= my_rom(9044); 
 data8 <= my_rom(10399); 
 data9 <= my_rom(11754); 
 data10 <= my_rom(13109);
when "01110010011" => 
 data1 <= my_rom(915); 
 data2 <= my_rom(2270); 
 data3 <= my_rom(3625); 
 data4 <= my_rom(4980); 
 data5 <= my_rom(6335); 
 data6 <= my_rom(7690); 
 data7 <= my_rom(9045); 
 data8 <= my_rom(10400); 
 data9 <= my_rom(11755); 
 data10 <= my_rom(13110);
when "01110010100" => 
 data1 <= my_rom(916); 
 data2 <= my_rom(2271); 
 data3 <= my_rom(3626); 
 data4 <= my_rom(4981); 
 data5 <= my_rom(6336); 
 data6 <= my_rom(7691); 
 data7 <= my_rom(9046); 
 data8 <= my_rom(10401); 
 data9 <= my_rom(11756); 
 data10 <= my_rom(13111);
when "01110010101" => 
 data1 <= my_rom(917); 
 data2 <= my_rom(2272); 
 data3 <= my_rom(3627); 
 data4 <= my_rom(4982); 
 data5 <= my_rom(6337); 
 data6 <= my_rom(7692); 
 data7 <= my_rom(9047); 
 data8 <= my_rom(10402); 
 data9 <= my_rom(11757); 
 data10 <= my_rom(13112);
when "01110010110" => 
 data1 <= my_rom(918); 
 data2 <= my_rom(2273); 
 data3 <= my_rom(3628); 
 data4 <= my_rom(4983); 
 data5 <= my_rom(6338); 
 data6 <= my_rom(7693); 
 data7 <= my_rom(9048); 
 data8 <= my_rom(10403); 
 data9 <= my_rom(11758); 
 data10 <= my_rom(13113);
when "01110010111" => 
 data1 <= my_rom(919); 
 data2 <= my_rom(2274); 
 data3 <= my_rom(3629); 
 data4 <= my_rom(4984); 
 data5 <= my_rom(6339); 
 data6 <= my_rom(7694); 
 data7 <= my_rom(9049); 
 data8 <= my_rom(10404); 
 data9 <= my_rom(11759); 
 data10 <= my_rom(13114);
when "01110011000" => 
 data1 <= my_rom(920); 
 data2 <= my_rom(2275); 
 data3 <= my_rom(3630); 
 data4 <= my_rom(4985); 
 data5 <= my_rom(6340); 
 data6 <= my_rom(7695); 
 data7 <= my_rom(9050); 
 data8 <= my_rom(10405); 
 data9 <= my_rom(11760); 
 data10 <= my_rom(13115);
when "01110011001" => 
 data1 <= my_rom(921); 
 data2 <= my_rom(2276); 
 data3 <= my_rom(3631); 
 data4 <= my_rom(4986); 
 data5 <= my_rom(6341); 
 data6 <= my_rom(7696); 
 data7 <= my_rom(9051); 
 data8 <= my_rom(10406); 
 data9 <= my_rom(11761); 
 data10 <= my_rom(13116);
when "01110011010" => 
 data1 <= my_rom(922); 
 data2 <= my_rom(2277); 
 data3 <= my_rom(3632); 
 data4 <= my_rom(4987); 
 data5 <= my_rom(6342); 
 data6 <= my_rom(7697); 
 data7 <= my_rom(9052); 
 data8 <= my_rom(10407); 
 data9 <= my_rom(11762); 
 data10 <= my_rom(13117);
when "01110011011" => 
 data1 <= my_rom(923); 
 data2 <= my_rom(2278); 
 data3 <= my_rom(3633); 
 data4 <= my_rom(4988); 
 data5 <= my_rom(6343); 
 data6 <= my_rom(7698); 
 data7 <= my_rom(9053); 
 data8 <= my_rom(10408); 
 data9 <= my_rom(11763); 
 data10 <= my_rom(13118);
when "01110011100" => 
 data1 <= my_rom(924); 
 data2 <= my_rom(2279); 
 data3 <= my_rom(3634); 
 data4 <= my_rom(4989); 
 data5 <= my_rom(6344); 
 data6 <= my_rom(7699); 
 data7 <= my_rom(9054); 
 data8 <= my_rom(10409); 
 data9 <= my_rom(11764); 
 data10 <= my_rom(13119);
when "01110011101" => 
 data1 <= my_rom(925); 
 data2 <= my_rom(2280); 
 data3 <= my_rom(3635); 
 data4 <= my_rom(4990); 
 data5 <= my_rom(6345); 
 data6 <= my_rom(7700); 
 data7 <= my_rom(9055); 
 data8 <= my_rom(10410); 
 data9 <= my_rom(11765); 
 data10 <= my_rom(13120);
when "01110011110" => 
 data1 <= my_rom(926); 
 data2 <= my_rom(2281); 
 data3 <= my_rom(3636); 
 data4 <= my_rom(4991); 
 data5 <= my_rom(6346); 
 data6 <= my_rom(7701); 
 data7 <= my_rom(9056); 
 data8 <= my_rom(10411); 
 data9 <= my_rom(11766); 
 data10 <= my_rom(13121);
when "01110011111" => 
 data1 <= my_rom(927); 
 data2 <= my_rom(2282); 
 data3 <= my_rom(3637); 
 data4 <= my_rom(4992); 
 data5 <= my_rom(6347); 
 data6 <= my_rom(7702); 
 data7 <= my_rom(9057); 
 data8 <= my_rom(10412); 
 data9 <= my_rom(11767); 
 data10 <= my_rom(13122);
when "01110100000" => 
 data1 <= my_rom(928); 
 data2 <= my_rom(2283); 
 data3 <= my_rom(3638); 
 data4 <= my_rom(4993); 
 data5 <= my_rom(6348); 
 data6 <= my_rom(7703); 
 data7 <= my_rom(9058); 
 data8 <= my_rom(10413); 
 data9 <= my_rom(11768); 
 data10 <= my_rom(13123);
when "01110100001" => 
 data1 <= my_rom(929); 
 data2 <= my_rom(2284); 
 data3 <= my_rom(3639); 
 data4 <= my_rom(4994); 
 data5 <= my_rom(6349); 
 data6 <= my_rom(7704); 
 data7 <= my_rom(9059); 
 data8 <= my_rom(10414); 
 data9 <= my_rom(11769); 
 data10 <= my_rom(13124);
when "01110100010" => 
 data1 <= my_rom(930); 
 data2 <= my_rom(2285); 
 data3 <= my_rom(3640); 
 data4 <= my_rom(4995); 
 data5 <= my_rom(6350); 
 data6 <= my_rom(7705); 
 data7 <= my_rom(9060); 
 data8 <= my_rom(10415); 
 data9 <= my_rom(11770); 
 data10 <= my_rom(13125);
when "01110100011" => 
 data1 <= my_rom(931); 
 data2 <= my_rom(2286); 
 data3 <= my_rom(3641); 
 data4 <= my_rom(4996); 
 data5 <= my_rom(6351); 
 data6 <= my_rom(7706); 
 data7 <= my_rom(9061); 
 data8 <= my_rom(10416); 
 data9 <= my_rom(11771); 
 data10 <= my_rom(13126);
when "01110100100" => 
 data1 <= my_rom(932); 
 data2 <= my_rom(2287); 
 data3 <= my_rom(3642); 
 data4 <= my_rom(4997); 
 data5 <= my_rom(6352); 
 data6 <= my_rom(7707); 
 data7 <= my_rom(9062); 
 data8 <= my_rom(10417); 
 data9 <= my_rom(11772); 
 data10 <= my_rom(13127);
when "01110100101" => 
 data1 <= my_rom(933); 
 data2 <= my_rom(2288); 
 data3 <= my_rom(3643); 
 data4 <= my_rom(4998); 
 data5 <= my_rom(6353); 
 data6 <= my_rom(7708); 
 data7 <= my_rom(9063); 
 data8 <= my_rom(10418); 
 data9 <= my_rom(11773); 
 data10 <= my_rom(13128);
when "01110100110" => 
 data1 <= my_rom(934); 
 data2 <= my_rom(2289); 
 data3 <= my_rom(3644); 
 data4 <= my_rom(4999); 
 data5 <= my_rom(6354); 
 data6 <= my_rom(7709); 
 data7 <= my_rom(9064); 
 data8 <= my_rom(10419); 
 data9 <= my_rom(11774); 
 data10 <= my_rom(13129);
when "01110100111" => 
 data1 <= my_rom(935); 
 data2 <= my_rom(2290); 
 data3 <= my_rom(3645); 
 data4 <= my_rom(5000); 
 data5 <= my_rom(6355); 
 data6 <= my_rom(7710); 
 data7 <= my_rom(9065); 
 data8 <= my_rom(10420); 
 data9 <= my_rom(11775); 
 data10 <= my_rom(13130);
when "01110101000" => 
 data1 <= my_rom(936); 
 data2 <= my_rom(2291); 
 data3 <= my_rom(3646); 
 data4 <= my_rom(5001); 
 data5 <= my_rom(6356); 
 data6 <= my_rom(7711); 
 data7 <= my_rom(9066); 
 data8 <= my_rom(10421); 
 data9 <= my_rom(11776); 
 data10 <= my_rom(13131);
when "01110101001" => 
 data1 <= my_rom(937); 
 data2 <= my_rom(2292); 
 data3 <= my_rom(3647); 
 data4 <= my_rom(5002); 
 data5 <= my_rom(6357); 
 data6 <= my_rom(7712); 
 data7 <= my_rom(9067); 
 data8 <= my_rom(10422); 
 data9 <= my_rom(11777); 
 data10 <= my_rom(13132);
when "01110101010" => 
 data1 <= my_rom(938); 
 data2 <= my_rom(2293); 
 data3 <= my_rom(3648); 
 data4 <= my_rom(5003); 
 data5 <= my_rom(6358); 
 data6 <= my_rom(7713); 
 data7 <= my_rom(9068); 
 data8 <= my_rom(10423); 
 data9 <= my_rom(11778); 
 data10 <= my_rom(13133);
when "01110101011" => 
 data1 <= my_rom(939); 
 data2 <= my_rom(2294); 
 data3 <= my_rom(3649); 
 data4 <= my_rom(5004); 
 data5 <= my_rom(6359); 
 data6 <= my_rom(7714); 
 data7 <= my_rom(9069); 
 data8 <= my_rom(10424); 
 data9 <= my_rom(11779); 
 data10 <= my_rom(13134);
when "01110101100" => 
 data1 <= my_rom(940); 
 data2 <= my_rom(2295); 
 data3 <= my_rom(3650); 
 data4 <= my_rom(5005); 
 data5 <= my_rom(6360); 
 data6 <= my_rom(7715); 
 data7 <= my_rom(9070); 
 data8 <= my_rom(10425); 
 data9 <= my_rom(11780); 
 data10 <= my_rom(13135);
when "01110101101" => 
 data1 <= my_rom(941); 
 data2 <= my_rom(2296); 
 data3 <= my_rom(3651); 
 data4 <= my_rom(5006); 
 data5 <= my_rom(6361); 
 data6 <= my_rom(7716); 
 data7 <= my_rom(9071); 
 data8 <= my_rom(10426); 
 data9 <= my_rom(11781); 
 data10 <= my_rom(13136);
when "01110101110" => 
 data1 <= my_rom(942); 
 data2 <= my_rom(2297); 
 data3 <= my_rom(3652); 
 data4 <= my_rom(5007); 
 data5 <= my_rom(6362); 
 data6 <= my_rom(7717); 
 data7 <= my_rom(9072); 
 data8 <= my_rom(10427); 
 data9 <= my_rom(11782); 
 data10 <= my_rom(13137);
when "01110101111" => 
 data1 <= my_rom(943); 
 data2 <= my_rom(2298); 
 data3 <= my_rom(3653); 
 data4 <= my_rom(5008); 
 data5 <= my_rom(6363); 
 data6 <= my_rom(7718); 
 data7 <= my_rom(9073); 
 data8 <= my_rom(10428); 
 data9 <= my_rom(11783); 
 data10 <= my_rom(13138);
when "01110110000" => 
 data1 <= my_rom(944); 
 data2 <= my_rom(2299); 
 data3 <= my_rom(3654); 
 data4 <= my_rom(5009); 
 data5 <= my_rom(6364); 
 data6 <= my_rom(7719); 
 data7 <= my_rom(9074); 
 data8 <= my_rom(10429); 
 data9 <= my_rom(11784); 
 data10 <= my_rom(13139);
when "01110110001" => 
 data1 <= my_rom(945); 
 data2 <= my_rom(2300); 
 data3 <= my_rom(3655); 
 data4 <= my_rom(5010); 
 data5 <= my_rom(6365); 
 data6 <= my_rom(7720); 
 data7 <= my_rom(9075); 
 data8 <= my_rom(10430); 
 data9 <= my_rom(11785); 
 data10 <= my_rom(13140);
when "01110110010" => 
 data1 <= my_rom(946); 
 data2 <= my_rom(2301); 
 data3 <= my_rom(3656); 
 data4 <= my_rom(5011); 
 data5 <= my_rom(6366); 
 data6 <= my_rom(7721); 
 data7 <= my_rom(9076); 
 data8 <= my_rom(10431); 
 data9 <= my_rom(11786); 
 data10 <= my_rom(13141);
when "01110110011" => 
 data1 <= my_rom(947); 
 data2 <= my_rom(2302); 
 data3 <= my_rom(3657); 
 data4 <= my_rom(5012); 
 data5 <= my_rom(6367); 
 data6 <= my_rom(7722); 
 data7 <= my_rom(9077); 
 data8 <= my_rom(10432); 
 data9 <= my_rom(11787); 
 data10 <= my_rom(13142);
when "01110110100" => 
 data1 <= my_rom(948); 
 data2 <= my_rom(2303); 
 data3 <= my_rom(3658); 
 data4 <= my_rom(5013); 
 data5 <= my_rom(6368); 
 data6 <= my_rom(7723); 
 data7 <= my_rom(9078); 
 data8 <= my_rom(10433); 
 data9 <= my_rom(11788); 
 data10 <= my_rom(13143);
when "01110110101" => 
 data1 <= my_rom(949); 
 data2 <= my_rom(2304); 
 data3 <= my_rom(3659); 
 data4 <= my_rom(5014); 
 data5 <= my_rom(6369); 
 data6 <= my_rom(7724); 
 data7 <= my_rom(9079); 
 data8 <= my_rom(10434); 
 data9 <= my_rom(11789); 
 data10 <= my_rom(13144);
when "01110110110" => 
 data1 <= my_rom(950); 
 data2 <= my_rom(2305); 
 data3 <= my_rom(3660); 
 data4 <= my_rom(5015); 
 data5 <= my_rom(6370); 
 data6 <= my_rom(7725); 
 data7 <= my_rom(9080); 
 data8 <= my_rom(10435); 
 data9 <= my_rom(11790); 
 data10 <= my_rom(13145);
when "01110110111" => 
 data1 <= my_rom(951); 
 data2 <= my_rom(2306); 
 data3 <= my_rom(3661); 
 data4 <= my_rom(5016); 
 data5 <= my_rom(6371); 
 data6 <= my_rom(7726); 
 data7 <= my_rom(9081); 
 data8 <= my_rom(10436); 
 data9 <= my_rom(11791); 
 data10 <= my_rom(13146);
when "01110111000" => 
 data1 <= my_rom(952); 
 data2 <= my_rom(2307); 
 data3 <= my_rom(3662); 
 data4 <= my_rom(5017); 
 data5 <= my_rom(6372); 
 data6 <= my_rom(7727); 
 data7 <= my_rom(9082); 
 data8 <= my_rom(10437); 
 data9 <= my_rom(11792); 
 data10 <= my_rom(13147);
when "01110111001" => 
 data1 <= my_rom(953); 
 data2 <= my_rom(2308); 
 data3 <= my_rom(3663); 
 data4 <= my_rom(5018); 
 data5 <= my_rom(6373); 
 data6 <= my_rom(7728); 
 data7 <= my_rom(9083); 
 data8 <= my_rom(10438); 
 data9 <= my_rom(11793); 
 data10 <= my_rom(13148);
when "01110111010" => 
 data1 <= my_rom(954); 
 data2 <= my_rom(2309); 
 data3 <= my_rom(3664); 
 data4 <= my_rom(5019); 
 data5 <= my_rom(6374); 
 data6 <= my_rom(7729); 
 data7 <= my_rom(9084); 
 data8 <= my_rom(10439); 
 data9 <= my_rom(11794); 
 data10 <= my_rom(13149);
when "01110111011" => 
 data1 <= my_rom(955); 
 data2 <= my_rom(2310); 
 data3 <= my_rom(3665); 
 data4 <= my_rom(5020); 
 data5 <= my_rom(6375); 
 data6 <= my_rom(7730); 
 data7 <= my_rom(9085); 
 data8 <= my_rom(10440); 
 data9 <= my_rom(11795); 
 data10 <= my_rom(13150);
when "01110111100" => 
 data1 <= my_rom(956); 
 data2 <= my_rom(2311); 
 data3 <= my_rom(3666); 
 data4 <= my_rom(5021); 
 data5 <= my_rom(6376); 
 data6 <= my_rom(7731); 
 data7 <= my_rom(9086); 
 data8 <= my_rom(10441); 
 data9 <= my_rom(11796); 
 data10 <= my_rom(13151);
when "01110111101" => 
 data1 <= my_rom(957); 
 data2 <= my_rom(2312); 
 data3 <= my_rom(3667); 
 data4 <= my_rom(5022); 
 data5 <= my_rom(6377); 
 data6 <= my_rom(7732); 
 data7 <= my_rom(9087); 
 data8 <= my_rom(10442); 
 data9 <= my_rom(11797); 
 data10 <= my_rom(13152);
when "01110111110" => 
 data1 <= my_rom(958); 
 data2 <= my_rom(2313); 
 data3 <= my_rom(3668); 
 data4 <= my_rom(5023); 
 data5 <= my_rom(6378); 
 data6 <= my_rom(7733); 
 data7 <= my_rom(9088); 
 data8 <= my_rom(10443); 
 data9 <= my_rom(11798); 
 data10 <= my_rom(13153);
when "01110111111" => 
 data1 <= my_rom(959); 
 data2 <= my_rom(2314); 
 data3 <= my_rom(3669); 
 data4 <= my_rom(5024); 
 data5 <= my_rom(6379); 
 data6 <= my_rom(7734); 
 data7 <= my_rom(9089); 
 data8 <= my_rom(10444); 
 data9 <= my_rom(11799); 
 data10 <= my_rom(13154);
when "01111000000" => 
 data1 <= my_rom(960); 
 data2 <= my_rom(2315); 
 data3 <= my_rom(3670); 
 data4 <= my_rom(5025); 
 data5 <= my_rom(6380); 
 data6 <= my_rom(7735); 
 data7 <= my_rom(9090); 
 data8 <= my_rom(10445); 
 data9 <= my_rom(11800); 
 data10 <= my_rom(13155);
when "01111000001" => 
 data1 <= my_rom(961); 
 data2 <= my_rom(2316); 
 data3 <= my_rom(3671); 
 data4 <= my_rom(5026); 
 data5 <= my_rom(6381); 
 data6 <= my_rom(7736); 
 data7 <= my_rom(9091); 
 data8 <= my_rom(10446); 
 data9 <= my_rom(11801); 
 data10 <= my_rom(13156);
when "01111000010" => 
 data1 <= my_rom(962); 
 data2 <= my_rom(2317); 
 data3 <= my_rom(3672); 
 data4 <= my_rom(5027); 
 data5 <= my_rom(6382); 
 data6 <= my_rom(7737); 
 data7 <= my_rom(9092); 
 data8 <= my_rom(10447); 
 data9 <= my_rom(11802); 
 data10 <= my_rom(13157);
when "01111000011" => 
 data1 <= my_rom(963); 
 data2 <= my_rom(2318); 
 data3 <= my_rom(3673); 
 data4 <= my_rom(5028); 
 data5 <= my_rom(6383); 
 data6 <= my_rom(7738); 
 data7 <= my_rom(9093); 
 data8 <= my_rom(10448); 
 data9 <= my_rom(11803); 
 data10 <= my_rom(13158);
when "01111000100" => 
 data1 <= my_rom(964); 
 data2 <= my_rom(2319); 
 data3 <= my_rom(3674); 
 data4 <= my_rom(5029); 
 data5 <= my_rom(6384); 
 data6 <= my_rom(7739); 
 data7 <= my_rom(9094); 
 data8 <= my_rom(10449); 
 data9 <= my_rom(11804); 
 data10 <= my_rom(13159);
when "01111000101" => 
 data1 <= my_rom(965); 
 data2 <= my_rom(2320); 
 data3 <= my_rom(3675); 
 data4 <= my_rom(5030); 
 data5 <= my_rom(6385); 
 data6 <= my_rom(7740); 
 data7 <= my_rom(9095); 
 data8 <= my_rom(10450); 
 data9 <= my_rom(11805); 
 data10 <= my_rom(13160);
when "01111000110" => 
 data1 <= my_rom(966); 
 data2 <= my_rom(2321); 
 data3 <= my_rom(3676); 
 data4 <= my_rom(5031); 
 data5 <= my_rom(6386); 
 data6 <= my_rom(7741); 
 data7 <= my_rom(9096); 
 data8 <= my_rom(10451); 
 data9 <= my_rom(11806); 
 data10 <= my_rom(13161);
when "01111000111" => 
 data1 <= my_rom(967); 
 data2 <= my_rom(2322); 
 data3 <= my_rom(3677); 
 data4 <= my_rom(5032); 
 data5 <= my_rom(6387); 
 data6 <= my_rom(7742); 
 data7 <= my_rom(9097); 
 data8 <= my_rom(10452); 
 data9 <= my_rom(11807); 
 data10 <= my_rom(13162);
when "01111001000" => 
 data1 <= my_rom(968); 
 data2 <= my_rom(2323); 
 data3 <= my_rom(3678); 
 data4 <= my_rom(5033); 
 data5 <= my_rom(6388); 
 data6 <= my_rom(7743); 
 data7 <= my_rom(9098); 
 data8 <= my_rom(10453); 
 data9 <= my_rom(11808); 
 data10 <= my_rom(13163);
when "01111001001" => 
 data1 <= my_rom(969); 
 data2 <= my_rom(2324); 
 data3 <= my_rom(3679); 
 data4 <= my_rom(5034); 
 data5 <= my_rom(6389); 
 data6 <= my_rom(7744); 
 data7 <= my_rom(9099); 
 data8 <= my_rom(10454); 
 data9 <= my_rom(11809); 
 data10 <= my_rom(13164);
when "01111001010" => 
 data1 <= my_rom(970); 
 data2 <= my_rom(2325); 
 data3 <= my_rom(3680); 
 data4 <= my_rom(5035); 
 data5 <= my_rom(6390); 
 data6 <= my_rom(7745); 
 data7 <= my_rom(9100); 
 data8 <= my_rom(10455); 
 data9 <= my_rom(11810); 
 data10 <= my_rom(13165);
when "01111001011" => 
 data1 <= my_rom(971); 
 data2 <= my_rom(2326); 
 data3 <= my_rom(3681); 
 data4 <= my_rom(5036); 
 data5 <= my_rom(6391); 
 data6 <= my_rom(7746); 
 data7 <= my_rom(9101); 
 data8 <= my_rom(10456); 
 data9 <= my_rom(11811); 
 data10 <= my_rom(13166);
when "01111001100" => 
 data1 <= my_rom(972); 
 data2 <= my_rom(2327); 
 data3 <= my_rom(3682); 
 data4 <= my_rom(5037); 
 data5 <= my_rom(6392); 
 data6 <= my_rom(7747); 
 data7 <= my_rom(9102); 
 data8 <= my_rom(10457); 
 data9 <= my_rom(11812); 
 data10 <= my_rom(13167);
when "01111001101" => 
 data1 <= my_rom(973); 
 data2 <= my_rom(2328); 
 data3 <= my_rom(3683); 
 data4 <= my_rom(5038); 
 data5 <= my_rom(6393); 
 data6 <= my_rom(7748); 
 data7 <= my_rom(9103); 
 data8 <= my_rom(10458); 
 data9 <= my_rom(11813); 
 data10 <= my_rom(13168);
when "01111001110" => 
 data1 <= my_rom(974); 
 data2 <= my_rom(2329); 
 data3 <= my_rom(3684); 
 data4 <= my_rom(5039); 
 data5 <= my_rom(6394); 
 data6 <= my_rom(7749); 
 data7 <= my_rom(9104); 
 data8 <= my_rom(10459); 
 data9 <= my_rom(11814); 
 data10 <= my_rom(13169);
when "01111001111" => 
 data1 <= my_rom(975); 
 data2 <= my_rom(2330); 
 data3 <= my_rom(3685); 
 data4 <= my_rom(5040); 
 data5 <= my_rom(6395); 
 data6 <= my_rom(7750); 
 data7 <= my_rom(9105); 
 data8 <= my_rom(10460); 
 data9 <= my_rom(11815); 
 data10 <= my_rom(13170);
when "01111010000" => 
 data1 <= my_rom(976); 
 data2 <= my_rom(2331); 
 data3 <= my_rom(3686); 
 data4 <= my_rom(5041); 
 data5 <= my_rom(6396); 
 data6 <= my_rom(7751); 
 data7 <= my_rom(9106); 
 data8 <= my_rom(10461); 
 data9 <= my_rom(11816); 
 data10 <= my_rom(13171);
when "01111010001" => 
 data1 <= my_rom(977); 
 data2 <= my_rom(2332); 
 data3 <= my_rom(3687); 
 data4 <= my_rom(5042); 
 data5 <= my_rom(6397); 
 data6 <= my_rom(7752); 
 data7 <= my_rom(9107); 
 data8 <= my_rom(10462); 
 data9 <= my_rom(11817); 
 data10 <= my_rom(13172);
when "01111010010" => 
 data1 <= my_rom(978); 
 data2 <= my_rom(2333); 
 data3 <= my_rom(3688); 
 data4 <= my_rom(5043); 
 data5 <= my_rom(6398); 
 data6 <= my_rom(7753); 
 data7 <= my_rom(9108); 
 data8 <= my_rom(10463); 
 data9 <= my_rom(11818); 
 data10 <= my_rom(13173);
when "01111010011" => 
 data1 <= my_rom(979); 
 data2 <= my_rom(2334); 
 data3 <= my_rom(3689); 
 data4 <= my_rom(5044); 
 data5 <= my_rom(6399); 
 data6 <= my_rom(7754); 
 data7 <= my_rom(9109); 
 data8 <= my_rom(10464); 
 data9 <= my_rom(11819); 
 data10 <= my_rom(13174);
when "01111010100" => 
 data1 <= my_rom(980); 
 data2 <= my_rom(2335); 
 data3 <= my_rom(3690); 
 data4 <= my_rom(5045); 
 data5 <= my_rom(6400); 
 data6 <= my_rom(7755); 
 data7 <= my_rom(9110); 
 data8 <= my_rom(10465); 
 data9 <= my_rom(11820); 
 data10 <= my_rom(13175);
when "01111010101" => 
 data1 <= my_rom(981); 
 data2 <= my_rom(2336); 
 data3 <= my_rom(3691); 
 data4 <= my_rom(5046); 
 data5 <= my_rom(6401); 
 data6 <= my_rom(7756); 
 data7 <= my_rom(9111); 
 data8 <= my_rom(10466); 
 data9 <= my_rom(11821); 
 data10 <= my_rom(13176);
when "01111010110" => 
 data1 <= my_rom(982); 
 data2 <= my_rom(2337); 
 data3 <= my_rom(3692); 
 data4 <= my_rom(5047); 
 data5 <= my_rom(6402); 
 data6 <= my_rom(7757); 
 data7 <= my_rom(9112); 
 data8 <= my_rom(10467); 
 data9 <= my_rom(11822); 
 data10 <= my_rom(13177);
when "01111010111" => 
 data1 <= my_rom(983); 
 data2 <= my_rom(2338); 
 data3 <= my_rom(3693); 
 data4 <= my_rom(5048); 
 data5 <= my_rom(6403); 
 data6 <= my_rom(7758); 
 data7 <= my_rom(9113); 
 data8 <= my_rom(10468); 
 data9 <= my_rom(11823); 
 data10 <= my_rom(13178);
when "01111011000" => 
 data1 <= my_rom(984); 
 data2 <= my_rom(2339); 
 data3 <= my_rom(3694); 
 data4 <= my_rom(5049); 
 data5 <= my_rom(6404); 
 data6 <= my_rom(7759); 
 data7 <= my_rom(9114); 
 data8 <= my_rom(10469); 
 data9 <= my_rom(11824); 
 data10 <= my_rom(13179);
when "01111011001" => 
 data1 <= my_rom(985); 
 data2 <= my_rom(2340); 
 data3 <= my_rom(3695); 
 data4 <= my_rom(5050); 
 data5 <= my_rom(6405); 
 data6 <= my_rom(7760); 
 data7 <= my_rom(9115); 
 data8 <= my_rom(10470); 
 data9 <= my_rom(11825); 
 data10 <= my_rom(13180);
when "01111011010" => 
 data1 <= my_rom(986); 
 data2 <= my_rom(2341); 
 data3 <= my_rom(3696); 
 data4 <= my_rom(5051); 
 data5 <= my_rom(6406); 
 data6 <= my_rom(7761); 
 data7 <= my_rom(9116); 
 data8 <= my_rom(10471); 
 data9 <= my_rom(11826); 
 data10 <= my_rom(13181);
when "01111011011" => 
 data1 <= my_rom(987); 
 data2 <= my_rom(2342); 
 data3 <= my_rom(3697); 
 data4 <= my_rom(5052); 
 data5 <= my_rom(6407); 
 data6 <= my_rom(7762); 
 data7 <= my_rom(9117); 
 data8 <= my_rom(10472); 
 data9 <= my_rom(11827); 
 data10 <= my_rom(13182);
when "01111011100" => 
 data1 <= my_rom(988); 
 data2 <= my_rom(2343); 
 data3 <= my_rom(3698); 
 data4 <= my_rom(5053); 
 data5 <= my_rom(6408); 
 data6 <= my_rom(7763); 
 data7 <= my_rom(9118); 
 data8 <= my_rom(10473); 
 data9 <= my_rom(11828); 
 data10 <= my_rom(13183);
when "01111011101" => 
 data1 <= my_rom(989); 
 data2 <= my_rom(2344); 
 data3 <= my_rom(3699); 
 data4 <= my_rom(5054); 
 data5 <= my_rom(6409); 
 data6 <= my_rom(7764); 
 data7 <= my_rom(9119); 
 data8 <= my_rom(10474); 
 data9 <= my_rom(11829); 
 data10 <= my_rom(13184);
when "01111011110" => 
 data1 <= my_rom(990); 
 data2 <= my_rom(2345); 
 data3 <= my_rom(3700); 
 data4 <= my_rom(5055); 
 data5 <= my_rom(6410); 
 data6 <= my_rom(7765); 
 data7 <= my_rom(9120); 
 data8 <= my_rom(10475); 
 data9 <= my_rom(11830); 
 data10 <= my_rom(13185);
when "01111011111" => 
 data1 <= my_rom(991); 
 data2 <= my_rom(2346); 
 data3 <= my_rom(3701); 
 data4 <= my_rom(5056); 
 data5 <= my_rom(6411); 
 data6 <= my_rom(7766); 
 data7 <= my_rom(9121); 
 data8 <= my_rom(10476); 
 data9 <= my_rom(11831); 
 data10 <= my_rom(13186);
when "01111100000" => 
 data1 <= my_rom(992); 
 data2 <= my_rom(2347); 
 data3 <= my_rom(3702); 
 data4 <= my_rom(5057); 
 data5 <= my_rom(6412); 
 data6 <= my_rom(7767); 
 data7 <= my_rom(9122); 
 data8 <= my_rom(10477); 
 data9 <= my_rom(11832); 
 data10 <= my_rom(13187);
when "01111100001" => 
 data1 <= my_rom(993); 
 data2 <= my_rom(2348); 
 data3 <= my_rom(3703); 
 data4 <= my_rom(5058); 
 data5 <= my_rom(6413); 
 data6 <= my_rom(7768); 
 data7 <= my_rom(9123); 
 data8 <= my_rom(10478); 
 data9 <= my_rom(11833); 
 data10 <= my_rom(13188);
when "01111100010" => 
 data1 <= my_rom(994); 
 data2 <= my_rom(2349); 
 data3 <= my_rom(3704); 
 data4 <= my_rom(5059); 
 data5 <= my_rom(6414); 
 data6 <= my_rom(7769); 
 data7 <= my_rom(9124); 
 data8 <= my_rom(10479); 
 data9 <= my_rom(11834); 
 data10 <= my_rom(13189);
when "01111100011" => 
 data1 <= my_rom(995); 
 data2 <= my_rom(2350); 
 data3 <= my_rom(3705); 
 data4 <= my_rom(5060); 
 data5 <= my_rom(6415); 
 data6 <= my_rom(7770); 
 data7 <= my_rom(9125); 
 data8 <= my_rom(10480); 
 data9 <= my_rom(11835); 
 data10 <= my_rom(13190);
when "01111100100" => 
 data1 <= my_rom(996); 
 data2 <= my_rom(2351); 
 data3 <= my_rom(3706); 
 data4 <= my_rom(5061); 
 data5 <= my_rom(6416); 
 data6 <= my_rom(7771); 
 data7 <= my_rom(9126); 
 data8 <= my_rom(10481); 
 data9 <= my_rom(11836); 
 data10 <= my_rom(13191);
when "01111100101" => 
 data1 <= my_rom(997); 
 data2 <= my_rom(2352); 
 data3 <= my_rom(3707); 
 data4 <= my_rom(5062); 
 data5 <= my_rom(6417); 
 data6 <= my_rom(7772); 
 data7 <= my_rom(9127); 
 data8 <= my_rom(10482); 
 data9 <= my_rom(11837); 
 data10 <= my_rom(13192);
when "01111100110" => 
 data1 <= my_rom(998); 
 data2 <= my_rom(2353); 
 data3 <= my_rom(3708); 
 data4 <= my_rom(5063); 
 data5 <= my_rom(6418); 
 data6 <= my_rom(7773); 
 data7 <= my_rom(9128); 
 data8 <= my_rom(10483); 
 data9 <= my_rom(11838); 
 data10 <= my_rom(13193);
when "01111100111" => 
 data1 <= my_rom(999); 
 data2 <= my_rom(2354); 
 data3 <= my_rom(3709); 
 data4 <= my_rom(5064); 
 data5 <= my_rom(6419); 
 data6 <= my_rom(7774); 
 data7 <= my_rom(9129); 
 data8 <= my_rom(10484); 
 data9 <= my_rom(11839); 
 data10 <= my_rom(13194);
when "01111101000" => 
 data1 <= my_rom(1000); 
 data2 <= my_rom(2355); 
 data3 <= my_rom(3710); 
 data4 <= my_rom(5065); 
 data5 <= my_rom(6420); 
 data6 <= my_rom(7775); 
 data7 <= my_rom(9130); 
 data8 <= my_rom(10485); 
 data9 <= my_rom(11840); 
 data10 <= my_rom(13195);
when "01111101001" => 
 data1 <= my_rom(1001); 
 data2 <= my_rom(2356); 
 data3 <= my_rom(3711); 
 data4 <= my_rom(5066); 
 data5 <= my_rom(6421); 
 data6 <= my_rom(7776); 
 data7 <= my_rom(9131); 
 data8 <= my_rom(10486); 
 data9 <= my_rom(11841); 
 data10 <= my_rom(13196);
when "01111101010" => 
 data1 <= my_rom(1002); 
 data2 <= my_rom(2357); 
 data3 <= my_rom(3712); 
 data4 <= my_rom(5067); 
 data5 <= my_rom(6422); 
 data6 <= my_rom(7777); 
 data7 <= my_rom(9132); 
 data8 <= my_rom(10487); 
 data9 <= my_rom(11842); 
 data10 <= my_rom(13197);
when "01111101011" => 
 data1 <= my_rom(1003); 
 data2 <= my_rom(2358); 
 data3 <= my_rom(3713); 
 data4 <= my_rom(5068); 
 data5 <= my_rom(6423); 
 data6 <= my_rom(7778); 
 data7 <= my_rom(9133); 
 data8 <= my_rom(10488); 
 data9 <= my_rom(11843); 
 data10 <= my_rom(13198);
when "01111101100" => 
 data1 <= my_rom(1004); 
 data2 <= my_rom(2359); 
 data3 <= my_rom(3714); 
 data4 <= my_rom(5069); 
 data5 <= my_rom(6424); 
 data6 <= my_rom(7779); 
 data7 <= my_rom(9134); 
 data8 <= my_rom(10489); 
 data9 <= my_rom(11844); 
 data10 <= my_rom(13199);
when "01111101101" => 
 data1 <= my_rom(1005); 
 data2 <= my_rom(2360); 
 data3 <= my_rom(3715); 
 data4 <= my_rom(5070); 
 data5 <= my_rom(6425); 
 data6 <= my_rom(7780); 
 data7 <= my_rom(9135); 
 data8 <= my_rom(10490); 
 data9 <= my_rom(11845); 
 data10 <= my_rom(13200);
when "01111101110" => 
 data1 <= my_rom(1006); 
 data2 <= my_rom(2361); 
 data3 <= my_rom(3716); 
 data4 <= my_rom(5071); 
 data5 <= my_rom(6426); 
 data6 <= my_rom(7781); 
 data7 <= my_rom(9136); 
 data8 <= my_rom(10491); 
 data9 <= my_rom(11846); 
 data10 <= my_rom(13201);
when "01111101111" => 
 data1 <= my_rom(1007); 
 data2 <= my_rom(2362); 
 data3 <= my_rom(3717); 
 data4 <= my_rom(5072); 
 data5 <= my_rom(6427); 
 data6 <= my_rom(7782); 
 data7 <= my_rom(9137); 
 data8 <= my_rom(10492); 
 data9 <= my_rom(11847); 
 data10 <= my_rom(13202);
when "01111110000" => 
 data1 <= my_rom(1008); 
 data2 <= my_rom(2363); 
 data3 <= my_rom(3718); 
 data4 <= my_rom(5073); 
 data5 <= my_rom(6428); 
 data6 <= my_rom(7783); 
 data7 <= my_rom(9138); 
 data8 <= my_rom(10493); 
 data9 <= my_rom(11848); 
 data10 <= my_rom(13203);
when "01111110001" => 
 data1 <= my_rom(1009); 
 data2 <= my_rom(2364); 
 data3 <= my_rom(3719); 
 data4 <= my_rom(5074); 
 data5 <= my_rom(6429); 
 data6 <= my_rom(7784); 
 data7 <= my_rom(9139); 
 data8 <= my_rom(10494); 
 data9 <= my_rom(11849); 
 data10 <= my_rom(13204);
when "01111110010" => 
 data1 <= my_rom(1010); 
 data2 <= my_rom(2365); 
 data3 <= my_rom(3720); 
 data4 <= my_rom(5075); 
 data5 <= my_rom(6430); 
 data6 <= my_rom(7785); 
 data7 <= my_rom(9140); 
 data8 <= my_rom(10495); 
 data9 <= my_rom(11850); 
 data10 <= my_rom(13205);
when "01111110011" => 
 data1 <= my_rom(1011); 
 data2 <= my_rom(2366); 
 data3 <= my_rom(3721); 
 data4 <= my_rom(5076); 
 data5 <= my_rom(6431); 
 data6 <= my_rom(7786); 
 data7 <= my_rom(9141); 
 data8 <= my_rom(10496); 
 data9 <= my_rom(11851); 
 data10 <= my_rom(13206);
when "01111110100" => 
 data1 <= my_rom(1012); 
 data2 <= my_rom(2367); 
 data3 <= my_rom(3722); 
 data4 <= my_rom(5077); 
 data5 <= my_rom(6432); 
 data6 <= my_rom(7787); 
 data7 <= my_rom(9142); 
 data8 <= my_rom(10497); 
 data9 <= my_rom(11852); 
 data10 <= my_rom(13207);
when "01111110101" => 
 data1 <= my_rom(1013); 
 data2 <= my_rom(2368); 
 data3 <= my_rom(3723); 
 data4 <= my_rom(5078); 
 data5 <= my_rom(6433); 
 data6 <= my_rom(7788); 
 data7 <= my_rom(9143); 
 data8 <= my_rom(10498); 
 data9 <= my_rom(11853); 
 data10 <= my_rom(13208);
when "01111110110" => 
 data1 <= my_rom(1014); 
 data2 <= my_rom(2369); 
 data3 <= my_rom(3724); 
 data4 <= my_rom(5079); 
 data5 <= my_rom(6434); 
 data6 <= my_rom(7789); 
 data7 <= my_rom(9144); 
 data8 <= my_rom(10499); 
 data9 <= my_rom(11854); 
 data10 <= my_rom(13209);
when "01111110111" => 
 data1 <= my_rom(1015); 
 data2 <= my_rom(2370); 
 data3 <= my_rom(3725); 
 data4 <= my_rom(5080); 
 data5 <= my_rom(6435); 
 data6 <= my_rom(7790); 
 data7 <= my_rom(9145); 
 data8 <= my_rom(10500); 
 data9 <= my_rom(11855); 
 data10 <= my_rom(13210);
when "01111111000" => 
 data1 <= my_rom(1016); 
 data2 <= my_rom(2371); 
 data3 <= my_rom(3726); 
 data4 <= my_rom(5081); 
 data5 <= my_rom(6436); 
 data6 <= my_rom(7791); 
 data7 <= my_rom(9146); 
 data8 <= my_rom(10501); 
 data9 <= my_rom(11856); 
 data10 <= my_rom(13211);
when "01111111001" => 
 data1 <= my_rom(1017); 
 data2 <= my_rom(2372); 
 data3 <= my_rom(3727); 
 data4 <= my_rom(5082); 
 data5 <= my_rom(6437); 
 data6 <= my_rom(7792); 
 data7 <= my_rom(9147); 
 data8 <= my_rom(10502); 
 data9 <= my_rom(11857); 
 data10 <= my_rom(13212);
when "01111111010" => 
 data1 <= my_rom(1018); 
 data2 <= my_rom(2373); 
 data3 <= my_rom(3728); 
 data4 <= my_rom(5083); 
 data5 <= my_rom(6438); 
 data6 <= my_rom(7793); 
 data7 <= my_rom(9148); 
 data8 <= my_rom(10503); 
 data9 <= my_rom(11858); 
 data10 <= my_rom(13213);
when "01111111011" => 
 data1 <= my_rom(1019); 
 data2 <= my_rom(2374); 
 data3 <= my_rom(3729); 
 data4 <= my_rom(5084); 
 data5 <= my_rom(6439); 
 data6 <= my_rom(7794); 
 data7 <= my_rom(9149); 
 data8 <= my_rom(10504); 
 data9 <= my_rom(11859); 
 data10 <= my_rom(13214);
when "01111111100" => 
 data1 <= my_rom(1020); 
 data2 <= my_rom(2375); 
 data3 <= my_rom(3730); 
 data4 <= my_rom(5085); 
 data5 <= my_rom(6440); 
 data6 <= my_rom(7795); 
 data7 <= my_rom(9150); 
 data8 <= my_rom(10505); 
 data9 <= my_rom(11860); 
 data10 <= my_rom(13215);
when "01111111101" => 
 data1 <= my_rom(1021); 
 data2 <= my_rom(2376); 
 data3 <= my_rom(3731); 
 data4 <= my_rom(5086); 
 data5 <= my_rom(6441); 
 data6 <= my_rom(7796); 
 data7 <= my_rom(9151); 
 data8 <= my_rom(10506); 
 data9 <= my_rom(11861); 
 data10 <= my_rom(13216);
when "01111111110" => 
 data1 <= my_rom(1022); 
 data2 <= my_rom(2377); 
 data3 <= my_rom(3732); 
 data4 <= my_rom(5087); 
 data5 <= my_rom(6442); 
 data6 <= my_rom(7797); 
 data7 <= my_rom(9152); 
 data8 <= my_rom(10507); 
 data9 <= my_rom(11862); 
 data10 <= my_rom(13217);
when "01111111111" => 
 data1 <= my_rom(1023); 
 data2 <= my_rom(2378); 
 data3 <= my_rom(3733); 
 data4 <= my_rom(5088); 
 data5 <= my_rom(6443); 
 data6 <= my_rom(7798); 
 data7 <= my_rom(9153); 
 data8 <= my_rom(10508); 
 data9 <= my_rom(11863); 
 data10 <= my_rom(13218);
when "10000000000" => 
 data1 <= my_rom(1024); 
 data2 <= my_rom(2379); 
 data3 <= my_rom(3734); 
 data4 <= my_rom(5089); 
 data5 <= my_rom(6444); 
 data6 <= my_rom(7799); 
 data7 <= my_rom(9154); 
 data8 <= my_rom(10509); 
 data9 <= my_rom(11864); 
 data10 <= my_rom(13219);
when "10000000001" => 
 data1 <= my_rom(1025); 
 data2 <= my_rom(2380); 
 data3 <= my_rom(3735); 
 data4 <= my_rom(5090); 
 data5 <= my_rom(6445); 
 data6 <= my_rom(7800); 
 data7 <= my_rom(9155); 
 data8 <= my_rom(10510); 
 data9 <= my_rom(11865); 
 data10 <= my_rom(13220);
when "10000000010" => 
 data1 <= my_rom(1026); 
 data2 <= my_rom(2381); 
 data3 <= my_rom(3736); 
 data4 <= my_rom(5091); 
 data5 <= my_rom(6446); 
 data6 <= my_rom(7801); 
 data7 <= my_rom(9156); 
 data8 <= my_rom(10511); 
 data9 <= my_rom(11866); 
 data10 <= my_rom(13221);
when "10000000011" => 
 data1 <= my_rom(1027); 
 data2 <= my_rom(2382); 
 data3 <= my_rom(3737); 
 data4 <= my_rom(5092); 
 data5 <= my_rom(6447); 
 data6 <= my_rom(7802); 
 data7 <= my_rom(9157); 
 data8 <= my_rom(10512); 
 data9 <= my_rom(11867); 
 data10 <= my_rom(13222);
when "10000000100" => 
 data1 <= my_rom(1028); 
 data2 <= my_rom(2383); 
 data3 <= my_rom(3738); 
 data4 <= my_rom(5093); 
 data5 <= my_rom(6448); 
 data6 <= my_rom(7803); 
 data7 <= my_rom(9158); 
 data8 <= my_rom(10513); 
 data9 <= my_rom(11868); 
 data10 <= my_rom(13223);
when "10000000101" => 
 data1 <= my_rom(1029); 
 data2 <= my_rom(2384); 
 data3 <= my_rom(3739); 
 data4 <= my_rom(5094); 
 data5 <= my_rom(6449); 
 data6 <= my_rom(7804); 
 data7 <= my_rom(9159); 
 data8 <= my_rom(10514); 
 data9 <= my_rom(11869); 
 data10 <= my_rom(13224);
when "10000000110" => 
 data1 <= my_rom(1030); 
 data2 <= my_rom(2385); 
 data3 <= my_rom(3740); 
 data4 <= my_rom(5095); 
 data5 <= my_rom(6450); 
 data6 <= my_rom(7805); 
 data7 <= my_rom(9160); 
 data8 <= my_rom(10515); 
 data9 <= my_rom(11870); 
 data10 <= my_rom(13225);
when "10000000111" => 
 data1 <= my_rom(1031); 
 data2 <= my_rom(2386); 
 data3 <= my_rom(3741); 
 data4 <= my_rom(5096); 
 data5 <= my_rom(6451); 
 data6 <= my_rom(7806); 
 data7 <= my_rom(9161); 
 data8 <= my_rom(10516); 
 data9 <= my_rom(11871); 
 data10 <= my_rom(13226);
when "10000001000" => 
 data1 <= my_rom(1032); 
 data2 <= my_rom(2387); 
 data3 <= my_rom(3742); 
 data4 <= my_rom(5097); 
 data5 <= my_rom(6452); 
 data6 <= my_rom(7807); 
 data7 <= my_rom(9162); 
 data8 <= my_rom(10517); 
 data9 <= my_rom(11872); 
 data10 <= my_rom(13227);
when "10000001001" => 
 data1 <= my_rom(1033); 
 data2 <= my_rom(2388); 
 data3 <= my_rom(3743); 
 data4 <= my_rom(5098); 
 data5 <= my_rom(6453); 
 data6 <= my_rom(7808); 
 data7 <= my_rom(9163); 
 data8 <= my_rom(10518); 
 data9 <= my_rom(11873); 
 data10 <= my_rom(13228);
when "10000001010" => 
 data1 <= my_rom(1034); 
 data2 <= my_rom(2389); 
 data3 <= my_rom(3744); 
 data4 <= my_rom(5099); 
 data5 <= my_rom(6454); 
 data6 <= my_rom(7809); 
 data7 <= my_rom(9164); 
 data8 <= my_rom(10519); 
 data9 <= my_rom(11874); 
 data10 <= my_rom(13229);
when "10000001011" => 
 data1 <= my_rom(1035); 
 data2 <= my_rom(2390); 
 data3 <= my_rom(3745); 
 data4 <= my_rom(5100); 
 data5 <= my_rom(6455); 
 data6 <= my_rom(7810); 
 data7 <= my_rom(9165); 
 data8 <= my_rom(10520); 
 data9 <= my_rom(11875); 
 data10 <= my_rom(13230);
when "10000001100" => 
 data1 <= my_rom(1036); 
 data2 <= my_rom(2391); 
 data3 <= my_rom(3746); 
 data4 <= my_rom(5101); 
 data5 <= my_rom(6456); 
 data6 <= my_rom(7811); 
 data7 <= my_rom(9166); 
 data8 <= my_rom(10521); 
 data9 <= my_rom(11876); 
 data10 <= my_rom(13231);
when "10000001101" => 
 data1 <= my_rom(1037); 
 data2 <= my_rom(2392); 
 data3 <= my_rom(3747); 
 data4 <= my_rom(5102); 
 data5 <= my_rom(6457); 
 data6 <= my_rom(7812); 
 data7 <= my_rom(9167); 
 data8 <= my_rom(10522); 
 data9 <= my_rom(11877); 
 data10 <= my_rom(13232);
when "10000001110" => 
 data1 <= my_rom(1038); 
 data2 <= my_rom(2393); 
 data3 <= my_rom(3748); 
 data4 <= my_rom(5103); 
 data5 <= my_rom(6458); 
 data6 <= my_rom(7813); 
 data7 <= my_rom(9168); 
 data8 <= my_rom(10523); 
 data9 <= my_rom(11878); 
 data10 <= my_rom(13233);
when "10000001111" => 
 data1 <= my_rom(1039); 
 data2 <= my_rom(2394); 
 data3 <= my_rom(3749); 
 data4 <= my_rom(5104); 
 data5 <= my_rom(6459); 
 data6 <= my_rom(7814); 
 data7 <= my_rom(9169); 
 data8 <= my_rom(10524); 
 data9 <= my_rom(11879); 
 data10 <= my_rom(13234);
when "10000010000" => 
 data1 <= my_rom(1040); 
 data2 <= my_rom(2395); 
 data3 <= my_rom(3750); 
 data4 <= my_rom(5105); 
 data5 <= my_rom(6460); 
 data6 <= my_rom(7815); 
 data7 <= my_rom(9170); 
 data8 <= my_rom(10525); 
 data9 <= my_rom(11880); 
 data10 <= my_rom(13235);
when "10000010001" => 
 data1 <= my_rom(1041); 
 data2 <= my_rom(2396); 
 data3 <= my_rom(3751); 
 data4 <= my_rom(5106); 
 data5 <= my_rom(6461); 
 data6 <= my_rom(7816); 
 data7 <= my_rom(9171); 
 data8 <= my_rom(10526); 
 data9 <= my_rom(11881); 
 data10 <= my_rom(13236);
when "10000010010" => 
 data1 <= my_rom(1042); 
 data2 <= my_rom(2397); 
 data3 <= my_rom(3752); 
 data4 <= my_rom(5107); 
 data5 <= my_rom(6462); 
 data6 <= my_rom(7817); 
 data7 <= my_rom(9172); 
 data8 <= my_rom(10527); 
 data9 <= my_rom(11882); 
 data10 <= my_rom(13237);
when "10000010011" => 
 data1 <= my_rom(1043); 
 data2 <= my_rom(2398); 
 data3 <= my_rom(3753); 
 data4 <= my_rom(5108); 
 data5 <= my_rom(6463); 
 data6 <= my_rom(7818); 
 data7 <= my_rom(9173); 
 data8 <= my_rom(10528); 
 data9 <= my_rom(11883); 
 data10 <= my_rom(13238);
when "10000010100" => 
 data1 <= my_rom(1044); 
 data2 <= my_rom(2399); 
 data3 <= my_rom(3754); 
 data4 <= my_rom(5109); 
 data5 <= my_rom(6464); 
 data6 <= my_rom(7819); 
 data7 <= my_rom(9174); 
 data8 <= my_rom(10529); 
 data9 <= my_rom(11884); 
 data10 <= my_rom(13239);
when "10000010101" => 
 data1 <= my_rom(1045); 
 data2 <= my_rom(2400); 
 data3 <= my_rom(3755); 
 data4 <= my_rom(5110); 
 data5 <= my_rom(6465); 
 data6 <= my_rom(7820); 
 data7 <= my_rom(9175); 
 data8 <= my_rom(10530); 
 data9 <= my_rom(11885); 
 data10 <= my_rom(13240);
when "10000010110" => 
 data1 <= my_rom(1046); 
 data2 <= my_rom(2401); 
 data3 <= my_rom(3756); 
 data4 <= my_rom(5111); 
 data5 <= my_rom(6466); 
 data6 <= my_rom(7821); 
 data7 <= my_rom(9176); 
 data8 <= my_rom(10531); 
 data9 <= my_rom(11886); 
 data10 <= my_rom(13241);
when "10000010111" => 
 data1 <= my_rom(1047); 
 data2 <= my_rom(2402); 
 data3 <= my_rom(3757); 
 data4 <= my_rom(5112); 
 data5 <= my_rom(6467); 
 data6 <= my_rom(7822); 
 data7 <= my_rom(9177); 
 data8 <= my_rom(10532); 
 data9 <= my_rom(11887); 
 data10 <= my_rom(13242);
when "10000011000" => 
 data1 <= my_rom(1048); 
 data2 <= my_rom(2403); 
 data3 <= my_rom(3758); 
 data4 <= my_rom(5113); 
 data5 <= my_rom(6468); 
 data6 <= my_rom(7823); 
 data7 <= my_rom(9178); 
 data8 <= my_rom(10533); 
 data9 <= my_rom(11888); 
 data10 <= my_rom(13243);
when "10000011001" => 
 data1 <= my_rom(1049); 
 data2 <= my_rom(2404); 
 data3 <= my_rom(3759); 
 data4 <= my_rom(5114); 
 data5 <= my_rom(6469); 
 data6 <= my_rom(7824); 
 data7 <= my_rom(9179); 
 data8 <= my_rom(10534); 
 data9 <= my_rom(11889); 
 data10 <= my_rom(13244);
when "10000011010" => 
 data1 <= my_rom(1050); 
 data2 <= my_rom(2405); 
 data3 <= my_rom(3760); 
 data4 <= my_rom(5115); 
 data5 <= my_rom(6470); 
 data6 <= my_rom(7825); 
 data7 <= my_rom(9180); 
 data8 <= my_rom(10535); 
 data9 <= my_rom(11890); 
 data10 <= my_rom(13245);
when "10000011011" => 
 data1 <= my_rom(1051); 
 data2 <= my_rom(2406); 
 data3 <= my_rom(3761); 
 data4 <= my_rom(5116); 
 data5 <= my_rom(6471); 
 data6 <= my_rom(7826); 
 data7 <= my_rom(9181); 
 data8 <= my_rom(10536); 
 data9 <= my_rom(11891); 
 data10 <= my_rom(13246);
when "10000011100" => 
 data1 <= my_rom(1052); 
 data2 <= my_rom(2407); 
 data3 <= my_rom(3762); 
 data4 <= my_rom(5117); 
 data5 <= my_rom(6472); 
 data6 <= my_rom(7827); 
 data7 <= my_rom(9182); 
 data8 <= my_rom(10537); 
 data9 <= my_rom(11892); 
 data10 <= my_rom(13247);
when "10000011101" => 
 data1 <= my_rom(1053); 
 data2 <= my_rom(2408); 
 data3 <= my_rom(3763); 
 data4 <= my_rom(5118); 
 data5 <= my_rom(6473); 
 data6 <= my_rom(7828); 
 data7 <= my_rom(9183); 
 data8 <= my_rom(10538); 
 data9 <= my_rom(11893); 
 data10 <= my_rom(13248);
when "10000011110" => 
 data1 <= my_rom(1054); 
 data2 <= my_rom(2409); 
 data3 <= my_rom(3764); 
 data4 <= my_rom(5119); 
 data5 <= my_rom(6474); 
 data6 <= my_rom(7829); 
 data7 <= my_rom(9184); 
 data8 <= my_rom(10539); 
 data9 <= my_rom(11894); 
 data10 <= my_rom(13249);
when "10000011111" => 
 data1 <= my_rom(1055); 
 data2 <= my_rom(2410); 
 data3 <= my_rom(3765); 
 data4 <= my_rom(5120); 
 data5 <= my_rom(6475); 
 data6 <= my_rom(7830); 
 data7 <= my_rom(9185); 
 data8 <= my_rom(10540); 
 data9 <= my_rom(11895); 
 data10 <= my_rom(13250);
when "10000100000" => 
 data1 <= my_rom(1056); 
 data2 <= my_rom(2411); 
 data3 <= my_rom(3766); 
 data4 <= my_rom(5121); 
 data5 <= my_rom(6476); 
 data6 <= my_rom(7831); 
 data7 <= my_rom(9186); 
 data8 <= my_rom(10541); 
 data9 <= my_rom(11896); 
 data10 <= my_rom(13251);
when "10000100001" => 
 data1 <= my_rom(1057); 
 data2 <= my_rom(2412); 
 data3 <= my_rom(3767); 
 data4 <= my_rom(5122); 
 data5 <= my_rom(6477); 
 data6 <= my_rom(7832); 
 data7 <= my_rom(9187); 
 data8 <= my_rom(10542); 
 data9 <= my_rom(11897); 
 data10 <= my_rom(13252);
when "10000100010" => 
 data1 <= my_rom(1058); 
 data2 <= my_rom(2413); 
 data3 <= my_rom(3768); 
 data4 <= my_rom(5123); 
 data5 <= my_rom(6478); 
 data6 <= my_rom(7833); 
 data7 <= my_rom(9188); 
 data8 <= my_rom(10543); 
 data9 <= my_rom(11898); 
 data10 <= my_rom(13253);
when "10000100011" => 
 data1 <= my_rom(1059); 
 data2 <= my_rom(2414); 
 data3 <= my_rom(3769); 
 data4 <= my_rom(5124); 
 data5 <= my_rom(6479); 
 data6 <= my_rom(7834); 
 data7 <= my_rom(9189); 
 data8 <= my_rom(10544); 
 data9 <= my_rom(11899); 
 data10 <= my_rom(13254);
when "10000100100" => 
 data1 <= my_rom(1060); 
 data2 <= my_rom(2415); 
 data3 <= my_rom(3770); 
 data4 <= my_rom(5125); 
 data5 <= my_rom(6480); 
 data6 <= my_rom(7835); 
 data7 <= my_rom(9190); 
 data8 <= my_rom(10545); 
 data9 <= my_rom(11900); 
 data10 <= my_rom(13255);
when "10000100101" => 
 data1 <= my_rom(1061); 
 data2 <= my_rom(2416); 
 data3 <= my_rom(3771); 
 data4 <= my_rom(5126); 
 data5 <= my_rom(6481); 
 data6 <= my_rom(7836); 
 data7 <= my_rom(9191); 
 data8 <= my_rom(10546); 
 data9 <= my_rom(11901); 
 data10 <= my_rom(13256);
when "10000100110" => 
 data1 <= my_rom(1062); 
 data2 <= my_rom(2417); 
 data3 <= my_rom(3772); 
 data4 <= my_rom(5127); 
 data5 <= my_rom(6482); 
 data6 <= my_rom(7837); 
 data7 <= my_rom(9192); 
 data8 <= my_rom(10547); 
 data9 <= my_rom(11902); 
 data10 <= my_rom(13257);
when "10000100111" => 
 data1 <= my_rom(1063); 
 data2 <= my_rom(2418); 
 data3 <= my_rom(3773); 
 data4 <= my_rom(5128); 
 data5 <= my_rom(6483); 
 data6 <= my_rom(7838); 
 data7 <= my_rom(9193); 
 data8 <= my_rom(10548); 
 data9 <= my_rom(11903); 
 data10 <= my_rom(13258);
when "10000101000" => 
 data1 <= my_rom(1064); 
 data2 <= my_rom(2419); 
 data3 <= my_rom(3774); 
 data4 <= my_rom(5129); 
 data5 <= my_rom(6484); 
 data6 <= my_rom(7839); 
 data7 <= my_rom(9194); 
 data8 <= my_rom(10549); 
 data9 <= my_rom(11904); 
 data10 <= my_rom(13259);
when "10000101001" => 
 data1 <= my_rom(1065); 
 data2 <= my_rom(2420); 
 data3 <= my_rom(3775); 
 data4 <= my_rom(5130); 
 data5 <= my_rom(6485); 
 data6 <= my_rom(7840); 
 data7 <= my_rom(9195); 
 data8 <= my_rom(10550); 
 data9 <= my_rom(11905); 
 data10 <= my_rom(13260);
when "10000101010" => 
 data1 <= my_rom(1066); 
 data2 <= my_rom(2421); 
 data3 <= my_rom(3776); 
 data4 <= my_rom(5131); 
 data5 <= my_rom(6486); 
 data6 <= my_rom(7841); 
 data7 <= my_rom(9196); 
 data8 <= my_rom(10551); 
 data9 <= my_rom(11906); 
 data10 <= my_rom(13261);
when "10000101011" => 
 data1 <= my_rom(1067); 
 data2 <= my_rom(2422); 
 data3 <= my_rom(3777); 
 data4 <= my_rom(5132); 
 data5 <= my_rom(6487); 
 data6 <= my_rom(7842); 
 data7 <= my_rom(9197); 
 data8 <= my_rom(10552); 
 data9 <= my_rom(11907); 
 data10 <= my_rom(13262);
when "10000101100" => 
 data1 <= my_rom(1068); 
 data2 <= my_rom(2423); 
 data3 <= my_rom(3778); 
 data4 <= my_rom(5133); 
 data5 <= my_rom(6488); 
 data6 <= my_rom(7843); 
 data7 <= my_rom(9198); 
 data8 <= my_rom(10553); 
 data9 <= my_rom(11908); 
 data10 <= my_rom(13263);
when "10000101101" => 
 data1 <= my_rom(1069); 
 data2 <= my_rom(2424); 
 data3 <= my_rom(3779); 
 data4 <= my_rom(5134); 
 data5 <= my_rom(6489); 
 data6 <= my_rom(7844); 
 data7 <= my_rom(9199); 
 data8 <= my_rom(10554); 
 data9 <= my_rom(11909); 
 data10 <= my_rom(13264);
when "10000101110" => 
 data1 <= my_rom(1070); 
 data2 <= my_rom(2425); 
 data3 <= my_rom(3780); 
 data4 <= my_rom(5135); 
 data5 <= my_rom(6490); 
 data6 <= my_rom(7845); 
 data7 <= my_rom(9200); 
 data8 <= my_rom(10555); 
 data9 <= my_rom(11910); 
 data10 <= my_rom(13265);
when "10000101111" => 
 data1 <= my_rom(1071); 
 data2 <= my_rom(2426); 
 data3 <= my_rom(3781); 
 data4 <= my_rom(5136); 
 data5 <= my_rom(6491); 
 data6 <= my_rom(7846); 
 data7 <= my_rom(9201); 
 data8 <= my_rom(10556); 
 data9 <= my_rom(11911); 
 data10 <= my_rom(13266);
when "10000110000" => 
 data1 <= my_rom(1072); 
 data2 <= my_rom(2427); 
 data3 <= my_rom(3782); 
 data4 <= my_rom(5137); 
 data5 <= my_rom(6492); 
 data6 <= my_rom(7847); 
 data7 <= my_rom(9202); 
 data8 <= my_rom(10557); 
 data9 <= my_rom(11912); 
 data10 <= my_rom(13267);
when "10000110001" => 
 data1 <= my_rom(1073); 
 data2 <= my_rom(2428); 
 data3 <= my_rom(3783); 
 data4 <= my_rom(5138); 
 data5 <= my_rom(6493); 
 data6 <= my_rom(7848); 
 data7 <= my_rom(9203); 
 data8 <= my_rom(10558); 
 data9 <= my_rom(11913); 
 data10 <= my_rom(13268);
when "10000110010" => 
 data1 <= my_rom(1074); 
 data2 <= my_rom(2429); 
 data3 <= my_rom(3784); 
 data4 <= my_rom(5139); 
 data5 <= my_rom(6494); 
 data6 <= my_rom(7849); 
 data7 <= my_rom(9204); 
 data8 <= my_rom(10559); 
 data9 <= my_rom(11914); 
 data10 <= my_rom(13269);
when "10000110011" => 
 data1 <= my_rom(1075); 
 data2 <= my_rom(2430); 
 data3 <= my_rom(3785); 
 data4 <= my_rom(5140); 
 data5 <= my_rom(6495); 
 data6 <= my_rom(7850); 
 data7 <= my_rom(9205); 
 data8 <= my_rom(10560); 
 data9 <= my_rom(11915); 
 data10 <= my_rom(13270);
when "10000110100" => 
 data1 <= my_rom(1076); 
 data2 <= my_rom(2431); 
 data3 <= my_rom(3786); 
 data4 <= my_rom(5141); 
 data5 <= my_rom(6496); 
 data6 <= my_rom(7851); 
 data7 <= my_rom(9206); 
 data8 <= my_rom(10561); 
 data9 <= my_rom(11916); 
 data10 <= my_rom(13271);
when "10000110101" => 
 data1 <= my_rom(1077); 
 data2 <= my_rom(2432); 
 data3 <= my_rom(3787); 
 data4 <= my_rom(5142); 
 data5 <= my_rom(6497); 
 data6 <= my_rom(7852); 
 data7 <= my_rom(9207); 
 data8 <= my_rom(10562); 
 data9 <= my_rom(11917); 
 data10 <= my_rom(13272);
when "10000110110" => 
 data1 <= my_rom(1078); 
 data2 <= my_rom(2433); 
 data3 <= my_rom(3788); 
 data4 <= my_rom(5143); 
 data5 <= my_rom(6498); 
 data6 <= my_rom(7853); 
 data7 <= my_rom(9208); 
 data8 <= my_rom(10563); 
 data9 <= my_rom(11918); 
 data10 <= my_rom(13273);
when "10000110111" => 
 data1 <= my_rom(1079); 
 data2 <= my_rom(2434); 
 data3 <= my_rom(3789); 
 data4 <= my_rom(5144); 
 data5 <= my_rom(6499); 
 data6 <= my_rom(7854); 
 data7 <= my_rom(9209); 
 data8 <= my_rom(10564); 
 data9 <= my_rom(11919); 
 data10 <= my_rom(13274);
when "10000111000" => 
 data1 <= my_rom(1080); 
 data2 <= my_rom(2435); 
 data3 <= my_rom(3790); 
 data4 <= my_rom(5145); 
 data5 <= my_rom(6500); 
 data6 <= my_rom(7855); 
 data7 <= my_rom(9210); 
 data8 <= my_rom(10565); 
 data9 <= my_rom(11920); 
 data10 <= my_rom(13275);
when "10000111001" => 
 data1 <= my_rom(1081); 
 data2 <= my_rom(2436); 
 data3 <= my_rom(3791); 
 data4 <= my_rom(5146); 
 data5 <= my_rom(6501); 
 data6 <= my_rom(7856); 
 data7 <= my_rom(9211); 
 data8 <= my_rom(10566); 
 data9 <= my_rom(11921); 
 data10 <= my_rom(13276);
when "10000111010" => 
 data1 <= my_rom(1082); 
 data2 <= my_rom(2437); 
 data3 <= my_rom(3792); 
 data4 <= my_rom(5147); 
 data5 <= my_rom(6502); 
 data6 <= my_rom(7857); 
 data7 <= my_rom(9212); 
 data8 <= my_rom(10567); 
 data9 <= my_rom(11922); 
 data10 <= my_rom(13277);
when "10000111011" => 
 data1 <= my_rom(1083); 
 data2 <= my_rom(2438); 
 data3 <= my_rom(3793); 
 data4 <= my_rom(5148); 
 data5 <= my_rom(6503); 
 data6 <= my_rom(7858); 
 data7 <= my_rom(9213); 
 data8 <= my_rom(10568); 
 data9 <= my_rom(11923); 
 data10 <= my_rom(13278);
when "10000111100" => 
 data1 <= my_rom(1084); 
 data2 <= my_rom(2439); 
 data3 <= my_rom(3794); 
 data4 <= my_rom(5149); 
 data5 <= my_rom(6504); 
 data6 <= my_rom(7859); 
 data7 <= my_rom(9214); 
 data8 <= my_rom(10569); 
 data9 <= my_rom(11924); 
 data10 <= my_rom(13279);
when "10000111101" => 
 data1 <= my_rom(1085); 
 data2 <= my_rom(2440); 
 data3 <= my_rom(3795); 
 data4 <= my_rom(5150); 
 data5 <= my_rom(6505); 
 data6 <= my_rom(7860); 
 data7 <= my_rom(9215); 
 data8 <= my_rom(10570); 
 data9 <= my_rom(11925); 
 data10 <= my_rom(13280);
when "10000111110" => 
 data1 <= my_rom(1086); 
 data2 <= my_rom(2441); 
 data3 <= my_rom(3796); 
 data4 <= my_rom(5151); 
 data5 <= my_rom(6506); 
 data6 <= my_rom(7861); 
 data7 <= my_rom(9216); 
 data8 <= my_rom(10571); 
 data9 <= my_rom(11926); 
 data10 <= my_rom(13281);
when "10000111111" => 
 data1 <= my_rom(1087); 
 data2 <= my_rom(2442); 
 data3 <= my_rom(3797); 
 data4 <= my_rom(5152); 
 data5 <= my_rom(6507); 
 data6 <= my_rom(7862); 
 data7 <= my_rom(9217); 
 data8 <= my_rom(10572); 
 data9 <= my_rom(11927); 
 data10 <= my_rom(13282);
when "10001000000" => 
 data1 <= my_rom(1088); 
 data2 <= my_rom(2443); 
 data3 <= my_rom(3798); 
 data4 <= my_rom(5153); 
 data5 <= my_rom(6508); 
 data6 <= my_rom(7863); 
 data7 <= my_rom(9218); 
 data8 <= my_rom(10573); 
 data9 <= my_rom(11928); 
 data10 <= my_rom(13283);
when "10001000001" => 
 data1 <= my_rom(1089); 
 data2 <= my_rom(2444); 
 data3 <= my_rom(3799); 
 data4 <= my_rom(5154); 
 data5 <= my_rom(6509); 
 data6 <= my_rom(7864); 
 data7 <= my_rom(9219); 
 data8 <= my_rom(10574); 
 data9 <= my_rom(11929); 
 data10 <= my_rom(13284);
when "10001000010" => 
 data1 <= my_rom(1090); 
 data2 <= my_rom(2445); 
 data3 <= my_rom(3800); 
 data4 <= my_rom(5155); 
 data5 <= my_rom(6510); 
 data6 <= my_rom(7865); 
 data7 <= my_rom(9220); 
 data8 <= my_rom(10575); 
 data9 <= my_rom(11930); 
 data10 <= my_rom(13285);
when "10001000011" => 
 data1 <= my_rom(1091); 
 data2 <= my_rom(2446); 
 data3 <= my_rom(3801); 
 data4 <= my_rom(5156); 
 data5 <= my_rom(6511); 
 data6 <= my_rom(7866); 
 data7 <= my_rom(9221); 
 data8 <= my_rom(10576); 
 data9 <= my_rom(11931); 
 data10 <= my_rom(13286);
when "10001000100" => 
 data1 <= my_rom(1092); 
 data2 <= my_rom(2447); 
 data3 <= my_rom(3802); 
 data4 <= my_rom(5157); 
 data5 <= my_rom(6512); 
 data6 <= my_rom(7867); 
 data7 <= my_rom(9222); 
 data8 <= my_rom(10577); 
 data9 <= my_rom(11932); 
 data10 <= my_rom(13287);
when "10001000101" => 
 data1 <= my_rom(1093); 
 data2 <= my_rom(2448); 
 data3 <= my_rom(3803); 
 data4 <= my_rom(5158); 
 data5 <= my_rom(6513); 
 data6 <= my_rom(7868); 
 data7 <= my_rom(9223); 
 data8 <= my_rom(10578); 
 data9 <= my_rom(11933); 
 data10 <= my_rom(13288);
when "10001000110" => 
 data1 <= my_rom(1094); 
 data2 <= my_rom(2449); 
 data3 <= my_rom(3804); 
 data4 <= my_rom(5159); 
 data5 <= my_rom(6514); 
 data6 <= my_rom(7869); 
 data7 <= my_rom(9224); 
 data8 <= my_rom(10579); 
 data9 <= my_rom(11934); 
 data10 <= my_rom(13289);
when "10001000111" => 
 data1 <= my_rom(1095); 
 data2 <= my_rom(2450); 
 data3 <= my_rom(3805); 
 data4 <= my_rom(5160); 
 data5 <= my_rom(6515); 
 data6 <= my_rom(7870); 
 data7 <= my_rom(9225); 
 data8 <= my_rom(10580); 
 data9 <= my_rom(11935); 
 data10 <= my_rom(13290);
when "10001001000" => 
 data1 <= my_rom(1096); 
 data2 <= my_rom(2451); 
 data3 <= my_rom(3806); 
 data4 <= my_rom(5161); 
 data5 <= my_rom(6516); 
 data6 <= my_rom(7871); 
 data7 <= my_rom(9226); 
 data8 <= my_rom(10581); 
 data9 <= my_rom(11936); 
 data10 <= my_rom(13291);
when "10001001001" => 
 data1 <= my_rom(1097); 
 data2 <= my_rom(2452); 
 data3 <= my_rom(3807); 
 data4 <= my_rom(5162); 
 data5 <= my_rom(6517); 
 data6 <= my_rom(7872); 
 data7 <= my_rom(9227); 
 data8 <= my_rom(10582); 
 data9 <= my_rom(11937); 
 data10 <= my_rom(13292);
when "10001001010" => 
 data1 <= my_rom(1098); 
 data2 <= my_rom(2453); 
 data3 <= my_rom(3808); 
 data4 <= my_rom(5163); 
 data5 <= my_rom(6518); 
 data6 <= my_rom(7873); 
 data7 <= my_rom(9228); 
 data8 <= my_rom(10583); 
 data9 <= my_rom(11938); 
 data10 <= my_rom(13293);
when "10001001011" => 
 data1 <= my_rom(1099); 
 data2 <= my_rom(2454); 
 data3 <= my_rom(3809); 
 data4 <= my_rom(5164); 
 data5 <= my_rom(6519); 
 data6 <= my_rom(7874); 
 data7 <= my_rom(9229); 
 data8 <= my_rom(10584); 
 data9 <= my_rom(11939); 
 data10 <= my_rom(13294);
when "10001001100" => 
 data1 <= my_rom(1100); 
 data2 <= my_rom(2455); 
 data3 <= my_rom(3810); 
 data4 <= my_rom(5165); 
 data5 <= my_rom(6520); 
 data6 <= my_rom(7875); 
 data7 <= my_rom(9230); 
 data8 <= my_rom(10585); 
 data9 <= my_rom(11940); 
 data10 <= my_rom(13295);
when "10001001101" => 
 data1 <= my_rom(1101); 
 data2 <= my_rom(2456); 
 data3 <= my_rom(3811); 
 data4 <= my_rom(5166); 
 data5 <= my_rom(6521); 
 data6 <= my_rom(7876); 
 data7 <= my_rom(9231); 
 data8 <= my_rom(10586); 
 data9 <= my_rom(11941); 
 data10 <= my_rom(13296);
when "10001001110" => 
 data1 <= my_rom(1102); 
 data2 <= my_rom(2457); 
 data3 <= my_rom(3812); 
 data4 <= my_rom(5167); 
 data5 <= my_rom(6522); 
 data6 <= my_rom(7877); 
 data7 <= my_rom(9232); 
 data8 <= my_rom(10587); 
 data9 <= my_rom(11942); 
 data10 <= my_rom(13297);
when "10001001111" => 
 data1 <= my_rom(1103); 
 data2 <= my_rom(2458); 
 data3 <= my_rom(3813); 
 data4 <= my_rom(5168); 
 data5 <= my_rom(6523); 
 data6 <= my_rom(7878); 
 data7 <= my_rom(9233); 
 data8 <= my_rom(10588); 
 data9 <= my_rom(11943); 
 data10 <= my_rom(13298);
when "10001010000" => 
 data1 <= my_rom(1104); 
 data2 <= my_rom(2459); 
 data3 <= my_rom(3814); 
 data4 <= my_rom(5169); 
 data5 <= my_rom(6524); 
 data6 <= my_rom(7879); 
 data7 <= my_rom(9234); 
 data8 <= my_rom(10589); 
 data9 <= my_rom(11944); 
 data10 <= my_rom(13299);
when "10001010001" => 
 data1 <= my_rom(1105); 
 data2 <= my_rom(2460); 
 data3 <= my_rom(3815); 
 data4 <= my_rom(5170); 
 data5 <= my_rom(6525); 
 data6 <= my_rom(7880); 
 data7 <= my_rom(9235); 
 data8 <= my_rom(10590); 
 data9 <= my_rom(11945); 
 data10 <= my_rom(13300);
when "10001010010" => 
 data1 <= my_rom(1106); 
 data2 <= my_rom(2461); 
 data3 <= my_rom(3816); 
 data4 <= my_rom(5171); 
 data5 <= my_rom(6526); 
 data6 <= my_rom(7881); 
 data7 <= my_rom(9236); 
 data8 <= my_rom(10591); 
 data9 <= my_rom(11946); 
 data10 <= my_rom(13301);
when "10001010011" => 
 data1 <= my_rom(1107); 
 data2 <= my_rom(2462); 
 data3 <= my_rom(3817); 
 data4 <= my_rom(5172); 
 data5 <= my_rom(6527); 
 data6 <= my_rom(7882); 
 data7 <= my_rom(9237); 
 data8 <= my_rom(10592); 
 data9 <= my_rom(11947); 
 data10 <= my_rom(13302);
when "10001010100" => 
 data1 <= my_rom(1108); 
 data2 <= my_rom(2463); 
 data3 <= my_rom(3818); 
 data4 <= my_rom(5173); 
 data5 <= my_rom(6528); 
 data6 <= my_rom(7883); 
 data7 <= my_rom(9238); 
 data8 <= my_rom(10593); 
 data9 <= my_rom(11948); 
 data10 <= my_rom(13303);
when "10001010101" => 
 data1 <= my_rom(1109); 
 data2 <= my_rom(2464); 
 data3 <= my_rom(3819); 
 data4 <= my_rom(5174); 
 data5 <= my_rom(6529); 
 data6 <= my_rom(7884); 
 data7 <= my_rom(9239); 
 data8 <= my_rom(10594); 
 data9 <= my_rom(11949); 
 data10 <= my_rom(13304);
when "10001010110" => 
 data1 <= my_rom(1110); 
 data2 <= my_rom(2465); 
 data3 <= my_rom(3820); 
 data4 <= my_rom(5175); 
 data5 <= my_rom(6530); 
 data6 <= my_rom(7885); 
 data7 <= my_rom(9240); 
 data8 <= my_rom(10595); 
 data9 <= my_rom(11950); 
 data10 <= my_rom(13305);
when "10001010111" => 
 data1 <= my_rom(1111); 
 data2 <= my_rom(2466); 
 data3 <= my_rom(3821); 
 data4 <= my_rom(5176); 
 data5 <= my_rom(6531); 
 data6 <= my_rom(7886); 
 data7 <= my_rom(9241); 
 data8 <= my_rom(10596); 
 data9 <= my_rom(11951); 
 data10 <= my_rom(13306);
when "10001011000" => 
 data1 <= my_rom(1112); 
 data2 <= my_rom(2467); 
 data3 <= my_rom(3822); 
 data4 <= my_rom(5177); 
 data5 <= my_rom(6532); 
 data6 <= my_rom(7887); 
 data7 <= my_rom(9242); 
 data8 <= my_rom(10597); 
 data9 <= my_rom(11952); 
 data10 <= my_rom(13307);
when "10001011001" => 
 data1 <= my_rom(1113); 
 data2 <= my_rom(2468); 
 data3 <= my_rom(3823); 
 data4 <= my_rom(5178); 
 data5 <= my_rom(6533); 
 data6 <= my_rom(7888); 
 data7 <= my_rom(9243); 
 data8 <= my_rom(10598); 
 data9 <= my_rom(11953); 
 data10 <= my_rom(13308);
when "10001011010" => 
 data1 <= my_rom(1114); 
 data2 <= my_rom(2469); 
 data3 <= my_rom(3824); 
 data4 <= my_rom(5179); 
 data5 <= my_rom(6534); 
 data6 <= my_rom(7889); 
 data7 <= my_rom(9244); 
 data8 <= my_rom(10599); 
 data9 <= my_rom(11954); 
 data10 <= my_rom(13309);
when "10001011011" => 
 data1 <= my_rom(1115); 
 data2 <= my_rom(2470); 
 data3 <= my_rom(3825); 
 data4 <= my_rom(5180); 
 data5 <= my_rom(6535); 
 data6 <= my_rom(7890); 
 data7 <= my_rom(9245); 
 data8 <= my_rom(10600); 
 data9 <= my_rom(11955); 
 data10 <= my_rom(13310);
when "10001011100" => 
 data1 <= my_rom(1116); 
 data2 <= my_rom(2471); 
 data3 <= my_rom(3826); 
 data4 <= my_rom(5181); 
 data5 <= my_rom(6536); 
 data6 <= my_rom(7891); 
 data7 <= my_rom(9246); 
 data8 <= my_rom(10601); 
 data9 <= my_rom(11956); 
 data10 <= my_rom(13311);
when "10001011101" => 
 data1 <= my_rom(1117); 
 data2 <= my_rom(2472); 
 data3 <= my_rom(3827); 
 data4 <= my_rom(5182); 
 data5 <= my_rom(6537); 
 data6 <= my_rom(7892); 
 data7 <= my_rom(9247); 
 data8 <= my_rom(10602); 
 data9 <= my_rom(11957); 
 data10 <= my_rom(13312);
when "10001011110" => 
 data1 <= my_rom(1118); 
 data2 <= my_rom(2473); 
 data3 <= my_rom(3828); 
 data4 <= my_rom(5183); 
 data5 <= my_rom(6538); 
 data6 <= my_rom(7893); 
 data7 <= my_rom(9248); 
 data8 <= my_rom(10603); 
 data9 <= my_rom(11958); 
 data10 <= my_rom(13313);
when "10001011111" => 
 data1 <= my_rom(1119); 
 data2 <= my_rom(2474); 
 data3 <= my_rom(3829); 
 data4 <= my_rom(5184); 
 data5 <= my_rom(6539); 
 data6 <= my_rom(7894); 
 data7 <= my_rom(9249); 
 data8 <= my_rom(10604); 
 data9 <= my_rom(11959); 
 data10 <= my_rom(13314);
when "10001100000" => 
 data1 <= my_rom(1120); 
 data2 <= my_rom(2475); 
 data3 <= my_rom(3830); 
 data4 <= my_rom(5185); 
 data5 <= my_rom(6540); 
 data6 <= my_rom(7895); 
 data7 <= my_rom(9250); 
 data8 <= my_rom(10605); 
 data9 <= my_rom(11960); 
 data10 <= my_rom(13315);
when "10001100001" => 
 data1 <= my_rom(1121); 
 data2 <= my_rom(2476); 
 data3 <= my_rom(3831); 
 data4 <= my_rom(5186); 
 data5 <= my_rom(6541); 
 data6 <= my_rom(7896); 
 data7 <= my_rom(9251); 
 data8 <= my_rom(10606); 
 data9 <= my_rom(11961); 
 data10 <= my_rom(13316);
when "10001100010" => 
 data1 <= my_rom(1122); 
 data2 <= my_rom(2477); 
 data3 <= my_rom(3832); 
 data4 <= my_rom(5187); 
 data5 <= my_rom(6542); 
 data6 <= my_rom(7897); 
 data7 <= my_rom(9252); 
 data8 <= my_rom(10607); 
 data9 <= my_rom(11962); 
 data10 <= my_rom(13317);
when "10001100011" => 
 data1 <= my_rom(1123); 
 data2 <= my_rom(2478); 
 data3 <= my_rom(3833); 
 data4 <= my_rom(5188); 
 data5 <= my_rom(6543); 
 data6 <= my_rom(7898); 
 data7 <= my_rom(9253); 
 data8 <= my_rom(10608); 
 data9 <= my_rom(11963); 
 data10 <= my_rom(13318);
when "10001100100" => 
 data1 <= my_rom(1124); 
 data2 <= my_rom(2479); 
 data3 <= my_rom(3834); 
 data4 <= my_rom(5189); 
 data5 <= my_rom(6544); 
 data6 <= my_rom(7899); 
 data7 <= my_rom(9254); 
 data8 <= my_rom(10609); 
 data9 <= my_rom(11964); 
 data10 <= my_rom(13319);
when "10001100101" => 
 data1 <= my_rom(1125); 
 data2 <= my_rom(2480); 
 data3 <= my_rom(3835); 
 data4 <= my_rom(5190); 
 data5 <= my_rom(6545); 
 data6 <= my_rom(7900); 
 data7 <= my_rom(9255); 
 data8 <= my_rom(10610); 
 data9 <= my_rom(11965); 
 data10 <= my_rom(13320);
when "10001100110" => 
 data1 <= my_rom(1126); 
 data2 <= my_rom(2481); 
 data3 <= my_rom(3836); 
 data4 <= my_rom(5191); 
 data5 <= my_rom(6546); 
 data6 <= my_rom(7901); 
 data7 <= my_rom(9256); 
 data8 <= my_rom(10611); 
 data9 <= my_rom(11966); 
 data10 <= my_rom(13321);
when "10001100111" => 
 data1 <= my_rom(1127); 
 data2 <= my_rom(2482); 
 data3 <= my_rom(3837); 
 data4 <= my_rom(5192); 
 data5 <= my_rom(6547); 
 data6 <= my_rom(7902); 
 data7 <= my_rom(9257); 
 data8 <= my_rom(10612); 
 data9 <= my_rom(11967); 
 data10 <= my_rom(13322);
when "10001101000" => 
 data1 <= my_rom(1128); 
 data2 <= my_rom(2483); 
 data3 <= my_rom(3838); 
 data4 <= my_rom(5193); 
 data5 <= my_rom(6548); 
 data6 <= my_rom(7903); 
 data7 <= my_rom(9258); 
 data8 <= my_rom(10613); 
 data9 <= my_rom(11968); 
 data10 <= my_rom(13323);
when "10001101001" => 
 data1 <= my_rom(1129); 
 data2 <= my_rom(2484); 
 data3 <= my_rom(3839); 
 data4 <= my_rom(5194); 
 data5 <= my_rom(6549); 
 data6 <= my_rom(7904); 
 data7 <= my_rom(9259); 
 data8 <= my_rom(10614); 
 data9 <= my_rom(11969); 
 data10 <= my_rom(13324);
when "10001101010" => 
 data1 <= my_rom(1130); 
 data2 <= my_rom(2485); 
 data3 <= my_rom(3840); 
 data4 <= my_rom(5195); 
 data5 <= my_rom(6550); 
 data6 <= my_rom(7905); 
 data7 <= my_rom(9260); 
 data8 <= my_rom(10615); 
 data9 <= my_rom(11970); 
 data10 <= my_rom(13325);
when "10001101011" => 
 data1 <= my_rom(1131); 
 data2 <= my_rom(2486); 
 data3 <= my_rom(3841); 
 data4 <= my_rom(5196); 
 data5 <= my_rom(6551); 
 data6 <= my_rom(7906); 
 data7 <= my_rom(9261); 
 data8 <= my_rom(10616); 
 data9 <= my_rom(11971); 
 data10 <= my_rom(13326);
when "10001101100" => 
 data1 <= my_rom(1132); 
 data2 <= my_rom(2487); 
 data3 <= my_rom(3842); 
 data4 <= my_rom(5197); 
 data5 <= my_rom(6552); 
 data6 <= my_rom(7907); 
 data7 <= my_rom(9262); 
 data8 <= my_rom(10617); 
 data9 <= my_rom(11972); 
 data10 <= my_rom(13327);
when "10001101101" => 
 data1 <= my_rom(1133); 
 data2 <= my_rom(2488); 
 data3 <= my_rom(3843); 
 data4 <= my_rom(5198); 
 data5 <= my_rom(6553); 
 data6 <= my_rom(7908); 
 data7 <= my_rom(9263); 
 data8 <= my_rom(10618); 
 data9 <= my_rom(11973); 
 data10 <= my_rom(13328);
when "10001101110" => 
 data1 <= my_rom(1134); 
 data2 <= my_rom(2489); 
 data3 <= my_rom(3844); 
 data4 <= my_rom(5199); 
 data5 <= my_rom(6554); 
 data6 <= my_rom(7909); 
 data7 <= my_rom(9264); 
 data8 <= my_rom(10619); 
 data9 <= my_rom(11974); 
 data10 <= my_rom(13329);
when "10001101111" => 
 data1 <= my_rom(1135); 
 data2 <= my_rom(2490); 
 data3 <= my_rom(3845); 
 data4 <= my_rom(5200); 
 data5 <= my_rom(6555); 
 data6 <= my_rom(7910); 
 data7 <= my_rom(9265); 
 data8 <= my_rom(10620); 
 data9 <= my_rom(11975); 
 data10 <= my_rom(13330);
when "10001110000" => 
 data1 <= my_rom(1136); 
 data2 <= my_rom(2491); 
 data3 <= my_rom(3846); 
 data4 <= my_rom(5201); 
 data5 <= my_rom(6556); 
 data6 <= my_rom(7911); 
 data7 <= my_rom(9266); 
 data8 <= my_rom(10621); 
 data9 <= my_rom(11976); 
 data10 <= my_rom(13331);
when "10001110001" => 
 data1 <= my_rom(1137); 
 data2 <= my_rom(2492); 
 data3 <= my_rom(3847); 
 data4 <= my_rom(5202); 
 data5 <= my_rom(6557); 
 data6 <= my_rom(7912); 
 data7 <= my_rom(9267); 
 data8 <= my_rom(10622); 
 data9 <= my_rom(11977); 
 data10 <= my_rom(13332);
when "10001110010" => 
 data1 <= my_rom(1138); 
 data2 <= my_rom(2493); 
 data3 <= my_rom(3848); 
 data4 <= my_rom(5203); 
 data5 <= my_rom(6558); 
 data6 <= my_rom(7913); 
 data7 <= my_rom(9268); 
 data8 <= my_rom(10623); 
 data9 <= my_rom(11978); 
 data10 <= my_rom(13333);
when "10001110011" => 
 data1 <= my_rom(1139); 
 data2 <= my_rom(2494); 
 data3 <= my_rom(3849); 
 data4 <= my_rom(5204); 
 data5 <= my_rom(6559); 
 data6 <= my_rom(7914); 
 data7 <= my_rom(9269); 
 data8 <= my_rom(10624); 
 data9 <= my_rom(11979); 
 data10 <= my_rom(13334);
when "10001110100" => 
 data1 <= my_rom(1140); 
 data2 <= my_rom(2495); 
 data3 <= my_rom(3850); 
 data4 <= my_rom(5205); 
 data5 <= my_rom(6560); 
 data6 <= my_rom(7915); 
 data7 <= my_rom(9270); 
 data8 <= my_rom(10625); 
 data9 <= my_rom(11980); 
 data10 <= my_rom(13335);
when "10001110101" => 
 data1 <= my_rom(1141); 
 data2 <= my_rom(2496); 
 data3 <= my_rom(3851); 
 data4 <= my_rom(5206); 
 data5 <= my_rom(6561); 
 data6 <= my_rom(7916); 
 data7 <= my_rom(9271); 
 data8 <= my_rom(10626); 
 data9 <= my_rom(11981); 
 data10 <= my_rom(13336);
when "10001110110" => 
 data1 <= my_rom(1142); 
 data2 <= my_rom(2497); 
 data3 <= my_rom(3852); 
 data4 <= my_rom(5207); 
 data5 <= my_rom(6562); 
 data6 <= my_rom(7917); 
 data7 <= my_rom(9272); 
 data8 <= my_rom(10627); 
 data9 <= my_rom(11982); 
 data10 <= my_rom(13337);
when "10001110111" => 
 data1 <= my_rom(1143); 
 data2 <= my_rom(2498); 
 data3 <= my_rom(3853); 
 data4 <= my_rom(5208); 
 data5 <= my_rom(6563); 
 data6 <= my_rom(7918); 
 data7 <= my_rom(9273); 
 data8 <= my_rom(10628); 
 data9 <= my_rom(11983); 
 data10 <= my_rom(13338);
when "10001111000" => 
 data1 <= my_rom(1144); 
 data2 <= my_rom(2499); 
 data3 <= my_rom(3854); 
 data4 <= my_rom(5209); 
 data5 <= my_rom(6564); 
 data6 <= my_rom(7919); 
 data7 <= my_rom(9274); 
 data8 <= my_rom(10629); 
 data9 <= my_rom(11984); 
 data10 <= my_rom(13339);
when "10001111001" => 
 data1 <= my_rom(1145); 
 data2 <= my_rom(2500); 
 data3 <= my_rom(3855); 
 data4 <= my_rom(5210); 
 data5 <= my_rom(6565); 
 data6 <= my_rom(7920); 
 data7 <= my_rom(9275); 
 data8 <= my_rom(10630); 
 data9 <= my_rom(11985); 
 data10 <= my_rom(13340);
when "10001111010" => 
 data1 <= my_rom(1146); 
 data2 <= my_rom(2501); 
 data3 <= my_rom(3856); 
 data4 <= my_rom(5211); 
 data5 <= my_rom(6566); 
 data6 <= my_rom(7921); 
 data7 <= my_rom(9276); 
 data8 <= my_rom(10631); 
 data9 <= my_rom(11986); 
 data10 <= my_rom(13341);
when "10001111011" => 
 data1 <= my_rom(1147); 
 data2 <= my_rom(2502); 
 data3 <= my_rom(3857); 
 data4 <= my_rom(5212); 
 data5 <= my_rom(6567); 
 data6 <= my_rom(7922); 
 data7 <= my_rom(9277); 
 data8 <= my_rom(10632); 
 data9 <= my_rom(11987); 
 data10 <= my_rom(13342);
when "10001111100" => 
 data1 <= my_rom(1148); 
 data2 <= my_rom(2503); 
 data3 <= my_rom(3858); 
 data4 <= my_rom(5213); 
 data5 <= my_rom(6568); 
 data6 <= my_rom(7923); 
 data7 <= my_rom(9278); 
 data8 <= my_rom(10633); 
 data9 <= my_rom(11988); 
 data10 <= my_rom(13343);
when "10001111101" => 
 data1 <= my_rom(1149); 
 data2 <= my_rom(2504); 
 data3 <= my_rom(3859); 
 data4 <= my_rom(5214); 
 data5 <= my_rom(6569); 
 data6 <= my_rom(7924); 
 data7 <= my_rom(9279); 
 data8 <= my_rom(10634); 
 data9 <= my_rom(11989); 
 data10 <= my_rom(13344);
when "10001111110" => 
 data1 <= my_rom(1150); 
 data2 <= my_rom(2505); 
 data3 <= my_rom(3860); 
 data4 <= my_rom(5215); 
 data5 <= my_rom(6570); 
 data6 <= my_rom(7925); 
 data7 <= my_rom(9280); 
 data8 <= my_rom(10635); 
 data9 <= my_rom(11990); 
 data10 <= my_rom(13345);
when "10001111111" => 
 data1 <= my_rom(1151); 
 data2 <= my_rom(2506); 
 data3 <= my_rom(3861); 
 data4 <= my_rom(5216); 
 data5 <= my_rom(6571); 
 data6 <= my_rom(7926); 
 data7 <= my_rom(9281); 
 data8 <= my_rom(10636); 
 data9 <= my_rom(11991); 
 data10 <= my_rom(13346);
when "10010000000" => 
 data1 <= my_rom(1152); 
 data2 <= my_rom(2507); 
 data3 <= my_rom(3862); 
 data4 <= my_rom(5217); 
 data5 <= my_rom(6572); 
 data6 <= my_rom(7927); 
 data7 <= my_rom(9282); 
 data8 <= my_rom(10637); 
 data9 <= my_rom(11992); 
 data10 <= my_rom(13347);
when "10010000001" => 
 data1 <= my_rom(1153); 
 data2 <= my_rom(2508); 
 data3 <= my_rom(3863); 
 data4 <= my_rom(5218); 
 data5 <= my_rom(6573); 
 data6 <= my_rom(7928); 
 data7 <= my_rom(9283); 
 data8 <= my_rom(10638); 
 data9 <= my_rom(11993); 
 data10 <= my_rom(13348);
when "10010000010" => 
 data1 <= my_rom(1154); 
 data2 <= my_rom(2509); 
 data3 <= my_rom(3864); 
 data4 <= my_rom(5219); 
 data5 <= my_rom(6574); 
 data6 <= my_rom(7929); 
 data7 <= my_rom(9284); 
 data8 <= my_rom(10639); 
 data9 <= my_rom(11994); 
 data10 <= my_rom(13349);
when "10010000011" => 
 data1 <= my_rom(1155); 
 data2 <= my_rom(2510); 
 data3 <= my_rom(3865); 
 data4 <= my_rom(5220); 
 data5 <= my_rom(6575); 
 data6 <= my_rom(7930); 
 data7 <= my_rom(9285); 
 data8 <= my_rom(10640); 
 data9 <= my_rom(11995); 
 data10 <= my_rom(13350);
when "10010000100" => 
 data1 <= my_rom(1156); 
 data2 <= my_rom(2511); 
 data3 <= my_rom(3866); 
 data4 <= my_rom(5221); 
 data5 <= my_rom(6576); 
 data6 <= my_rom(7931); 
 data7 <= my_rom(9286); 
 data8 <= my_rom(10641); 
 data9 <= my_rom(11996); 
 data10 <= my_rom(13351);
when "10010000101" => 
 data1 <= my_rom(1157); 
 data2 <= my_rom(2512); 
 data3 <= my_rom(3867); 
 data4 <= my_rom(5222); 
 data5 <= my_rom(6577); 
 data6 <= my_rom(7932); 
 data7 <= my_rom(9287); 
 data8 <= my_rom(10642); 
 data9 <= my_rom(11997); 
 data10 <= my_rom(13352);
when "10010000110" => 
 data1 <= my_rom(1158); 
 data2 <= my_rom(2513); 
 data3 <= my_rom(3868); 
 data4 <= my_rom(5223); 
 data5 <= my_rom(6578); 
 data6 <= my_rom(7933); 
 data7 <= my_rom(9288); 
 data8 <= my_rom(10643); 
 data9 <= my_rom(11998); 
 data10 <= my_rom(13353);
when "10010000111" => 
 data1 <= my_rom(1159); 
 data2 <= my_rom(2514); 
 data3 <= my_rom(3869); 
 data4 <= my_rom(5224); 
 data5 <= my_rom(6579); 
 data6 <= my_rom(7934); 
 data7 <= my_rom(9289); 
 data8 <= my_rom(10644); 
 data9 <= my_rom(11999); 
 data10 <= my_rom(13354);
when "10010001000" => 
 data1 <= my_rom(1160); 
 data2 <= my_rom(2515); 
 data3 <= my_rom(3870); 
 data4 <= my_rom(5225); 
 data5 <= my_rom(6580); 
 data6 <= my_rom(7935); 
 data7 <= my_rom(9290); 
 data8 <= my_rom(10645); 
 data9 <= my_rom(12000); 
 data10 <= my_rom(13355);
when "10010001001" => 
 data1 <= my_rom(1161); 
 data2 <= my_rom(2516); 
 data3 <= my_rom(3871); 
 data4 <= my_rom(5226); 
 data5 <= my_rom(6581); 
 data6 <= my_rom(7936); 
 data7 <= my_rom(9291); 
 data8 <= my_rom(10646); 
 data9 <= my_rom(12001); 
 data10 <= my_rom(13356);
when "10010001010" => 
 data1 <= my_rom(1162); 
 data2 <= my_rom(2517); 
 data3 <= my_rom(3872); 
 data4 <= my_rom(5227); 
 data5 <= my_rom(6582); 
 data6 <= my_rom(7937); 
 data7 <= my_rom(9292); 
 data8 <= my_rom(10647); 
 data9 <= my_rom(12002); 
 data10 <= my_rom(13357);
when "10010001011" => 
 data1 <= my_rom(1163); 
 data2 <= my_rom(2518); 
 data3 <= my_rom(3873); 
 data4 <= my_rom(5228); 
 data5 <= my_rom(6583); 
 data6 <= my_rom(7938); 
 data7 <= my_rom(9293); 
 data8 <= my_rom(10648); 
 data9 <= my_rom(12003); 
 data10 <= my_rom(13358);
when "10010001100" => 
 data1 <= my_rom(1164); 
 data2 <= my_rom(2519); 
 data3 <= my_rom(3874); 
 data4 <= my_rom(5229); 
 data5 <= my_rom(6584); 
 data6 <= my_rom(7939); 
 data7 <= my_rom(9294); 
 data8 <= my_rom(10649); 
 data9 <= my_rom(12004); 
 data10 <= my_rom(13359);
when "10010001101" => 
 data1 <= my_rom(1165); 
 data2 <= my_rom(2520); 
 data3 <= my_rom(3875); 
 data4 <= my_rom(5230); 
 data5 <= my_rom(6585); 
 data6 <= my_rom(7940); 
 data7 <= my_rom(9295); 
 data8 <= my_rom(10650); 
 data9 <= my_rom(12005); 
 data10 <= my_rom(13360);
when "10010001110" => 
 data1 <= my_rom(1166); 
 data2 <= my_rom(2521); 
 data3 <= my_rom(3876); 
 data4 <= my_rom(5231); 
 data5 <= my_rom(6586); 
 data6 <= my_rom(7941); 
 data7 <= my_rom(9296); 
 data8 <= my_rom(10651); 
 data9 <= my_rom(12006); 
 data10 <= my_rom(13361);
when "10010001111" => 
 data1 <= my_rom(1167); 
 data2 <= my_rom(2522); 
 data3 <= my_rom(3877); 
 data4 <= my_rom(5232); 
 data5 <= my_rom(6587); 
 data6 <= my_rom(7942); 
 data7 <= my_rom(9297); 
 data8 <= my_rom(10652); 
 data9 <= my_rom(12007); 
 data10 <= my_rom(13362);
when "10010010000" => 
 data1 <= my_rom(1168); 
 data2 <= my_rom(2523); 
 data3 <= my_rom(3878); 
 data4 <= my_rom(5233); 
 data5 <= my_rom(6588); 
 data6 <= my_rom(7943); 
 data7 <= my_rom(9298); 
 data8 <= my_rom(10653); 
 data9 <= my_rom(12008); 
 data10 <= my_rom(13363);
when "10010010001" => 
 data1 <= my_rom(1169); 
 data2 <= my_rom(2524); 
 data3 <= my_rom(3879); 
 data4 <= my_rom(5234); 
 data5 <= my_rom(6589); 
 data6 <= my_rom(7944); 
 data7 <= my_rom(9299); 
 data8 <= my_rom(10654); 
 data9 <= my_rom(12009); 
 data10 <= my_rom(13364);
when "10010010010" => 
 data1 <= my_rom(1170); 
 data2 <= my_rom(2525); 
 data3 <= my_rom(3880); 
 data4 <= my_rom(5235); 
 data5 <= my_rom(6590); 
 data6 <= my_rom(7945); 
 data7 <= my_rom(9300); 
 data8 <= my_rom(10655); 
 data9 <= my_rom(12010); 
 data10 <= my_rom(13365);
when "10010010011" => 
 data1 <= my_rom(1171); 
 data2 <= my_rom(2526); 
 data3 <= my_rom(3881); 
 data4 <= my_rom(5236); 
 data5 <= my_rom(6591); 
 data6 <= my_rom(7946); 
 data7 <= my_rom(9301); 
 data8 <= my_rom(10656); 
 data9 <= my_rom(12011); 
 data10 <= my_rom(13366);
when "10010010100" => 
 data1 <= my_rom(1172); 
 data2 <= my_rom(2527); 
 data3 <= my_rom(3882); 
 data4 <= my_rom(5237); 
 data5 <= my_rom(6592); 
 data6 <= my_rom(7947); 
 data7 <= my_rom(9302); 
 data8 <= my_rom(10657); 
 data9 <= my_rom(12012); 
 data10 <= my_rom(13367);
when "10010010101" => 
 data1 <= my_rom(1173); 
 data2 <= my_rom(2528); 
 data3 <= my_rom(3883); 
 data4 <= my_rom(5238); 
 data5 <= my_rom(6593); 
 data6 <= my_rom(7948); 
 data7 <= my_rom(9303); 
 data8 <= my_rom(10658); 
 data9 <= my_rom(12013); 
 data10 <= my_rom(13368);
when "10010010110" => 
 data1 <= my_rom(1174); 
 data2 <= my_rom(2529); 
 data3 <= my_rom(3884); 
 data4 <= my_rom(5239); 
 data5 <= my_rom(6594); 
 data6 <= my_rom(7949); 
 data7 <= my_rom(9304); 
 data8 <= my_rom(10659); 
 data9 <= my_rom(12014); 
 data10 <= my_rom(13369);
when "10010010111" => 
 data1 <= my_rom(1175); 
 data2 <= my_rom(2530); 
 data3 <= my_rom(3885); 
 data4 <= my_rom(5240); 
 data5 <= my_rom(6595); 
 data6 <= my_rom(7950); 
 data7 <= my_rom(9305); 
 data8 <= my_rom(10660); 
 data9 <= my_rom(12015); 
 data10 <= my_rom(13370);
when "10010011000" => 
 data1 <= my_rom(1176); 
 data2 <= my_rom(2531); 
 data3 <= my_rom(3886); 
 data4 <= my_rom(5241); 
 data5 <= my_rom(6596); 
 data6 <= my_rom(7951); 
 data7 <= my_rom(9306); 
 data8 <= my_rom(10661); 
 data9 <= my_rom(12016); 
 data10 <= my_rom(13371);
when "10010011001" => 
 data1 <= my_rom(1177); 
 data2 <= my_rom(2532); 
 data3 <= my_rom(3887); 
 data4 <= my_rom(5242); 
 data5 <= my_rom(6597); 
 data6 <= my_rom(7952); 
 data7 <= my_rom(9307); 
 data8 <= my_rom(10662); 
 data9 <= my_rom(12017); 
 data10 <= my_rom(13372);
when "10010011010" => 
 data1 <= my_rom(1178); 
 data2 <= my_rom(2533); 
 data3 <= my_rom(3888); 
 data4 <= my_rom(5243); 
 data5 <= my_rom(6598); 
 data6 <= my_rom(7953); 
 data7 <= my_rom(9308); 
 data8 <= my_rom(10663); 
 data9 <= my_rom(12018); 
 data10 <= my_rom(13373);
when "10010011011" => 
 data1 <= my_rom(1179); 
 data2 <= my_rom(2534); 
 data3 <= my_rom(3889); 
 data4 <= my_rom(5244); 
 data5 <= my_rom(6599); 
 data6 <= my_rom(7954); 
 data7 <= my_rom(9309); 
 data8 <= my_rom(10664); 
 data9 <= my_rom(12019); 
 data10 <= my_rom(13374);
when "10010011100" => 
 data1 <= my_rom(1180); 
 data2 <= my_rom(2535); 
 data3 <= my_rom(3890); 
 data4 <= my_rom(5245); 
 data5 <= my_rom(6600); 
 data6 <= my_rom(7955); 
 data7 <= my_rom(9310); 
 data8 <= my_rom(10665); 
 data9 <= my_rom(12020); 
 data10 <= my_rom(13375);
when "10010011101" => 
 data1 <= my_rom(1181); 
 data2 <= my_rom(2536); 
 data3 <= my_rom(3891); 
 data4 <= my_rom(5246); 
 data5 <= my_rom(6601); 
 data6 <= my_rom(7956); 
 data7 <= my_rom(9311); 
 data8 <= my_rom(10666); 
 data9 <= my_rom(12021); 
 data10 <= my_rom(13376);
when "10010011110" => 
 data1 <= my_rom(1182); 
 data2 <= my_rom(2537); 
 data3 <= my_rom(3892); 
 data4 <= my_rom(5247); 
 data5 <= my_rom(6602); 
 data6 <= my_rom(7957); 
 data7 <= my_rom(9312); 
 data8 <= my_rom(10667); 
 data9 <= my_rom(12022); 
 data10 <= my_rom(13377);
when "10010011111" => 
 data1 <= my_rom(1183); 
 data2 <= my_rom(2538); 
 data3 <= my_rom(3893); 
 data4 <= my_rom(5248); 
 data5 <= my_rom(6603); 
 data6 <= my_rom(7958); 
 data7 <= my_rom(9313); 
 data8 <= my_rom(10668); 
 data9 <= my_rom(12023); 
 data10 <= my_rom(13378);
when "10010100000" => 
 data1 <= my_rom(1184); 
 data2 <= my_rom(2539); 
 data3 <= my_rom(3894); 
 data4 <= my_rom(5249); 
 data5 <= my_rom(6604); 
 data6 <= my_rom(7959); 
 data7 <= my_rom(9314); 
 data8 <= my_rom(10669); 
 data9 <= my_rom(12024); 
 data10 <= my_rom(13379);
when "10010100001" => 
 data1 <= my_rom(1185); 
 data2 <= my_rom(2540); 
 data3 <= my_rom(3895); 
 data4 <= my_rom(5250); 
 data5 <= my_rom(6605); 
 data6 <= my_rom(7960); 
 data7 <= my_rom(9315); 
 data8 <= my_rom(10670); 
 data9 <= my_rom(12025); 
 data10 <= my_rom(13380);
when "10010100010" => 
 data1 <= my_rom(1186); 
 data2 <= my_rom(2541); 
 data3 <= my_rom(3896); 
 data4 <= my_rom(5251); 
 data5 <= my_rom(6606); 
 data6 <= my_rom(7961); 
 data7 <= my_rom(9316); 
 data8 <= my_rom(10671); 
 data9 <= my_rom(12026); 
 data10 <= my_rom(13381);
when "10010100011" => 
 data1 <= my_rom(1187); 
 data2 <= my_rom(2542); 
 data3 <= my_rom(3897); 
 data4 <= my_rom(5252); 
 data5 <= my_rom(6607); 
 data6 <= my_rom(7962); 
 data7 <= my_rom(9317); 
 data8 <= my_rom(10672); 
 data9 <= my_rom(12027); 
 data10 <= my_rom(13382);
when "10010100100" => 
 data1 <= my_rom(1188); 
 data2 <= my_rom(2543); 
 data3 <= my_rom(3898); 
 data4 <= my_rom(5253); 
 data5 <= my_rom(6608); 
 data6 <= my_rom(7963); 
 data7 <= my_rom(9318); 
 data8 <= my_rom(10673); 
 data9 <= my_rom(12028); 
 data10 <= my_rom(13383);
when "10010100101" => 
 data1 <= my_rom(1189); 
 data2 <= my_rom(2544); 
 data3 <= my_rom(3899); 
 data4 <= my_rom(5254); 
 data5 <= my_rom(6609); 
 data6 <= my_rom(7964); 
 data7 <= my_rom(9319); 
 data8 <= my_rom(10674); 
 data9 <= my_rom(12029); 
 data10 <= my_rom(13384);
when "10010100110" => 
 data1 <= my_rom(1190); 
 data2 <= my_rom(2545); 
 data3 <= my_rom(3900); 
 data4 <= my_rom(5255); 
 data5 <= my_rom(6610); 
 data6 <= my_rom(7965); 
 data7 <= my_rom(9320); 
 data8 <= my_rom(10675); 
 data9 <= my_rom(12030); 
 data10 <= my_rom(13385);
when "10010100111" => 
 data1 <= my_rom(1191); 
 data2 <= my_rom(2546); 
 data3 <= my_rom(3901); 
 data4 <= my_rom(5256); 
 data5 <= my_rom(6611); 
 data6 <= my_rom(7966); 
 data7 <= my_rom(9321); 
 data8 <= my_rom(10676); 
 data9 <= my_rom(12031); 
 data10 <= my_rom(13386);
when "10010101000" => 
 data1 <= my_rom(1192); 
 data2 <= my_rom(2547); 
 data3 <= my_rom(3902); 
 data4 <= my_rom(5257); 
 data5 <= my_rom(6612); 
 data6 <= my_rom(7967); 
 data7 <= my_rom(9322); 
 data8 <= my_rom(10677); 
 data9 <= my_rom(12032); 
 data10 <= my_rom(13387);
when "10010101001" => 
 data1 <= my_rom(1193); 
 data2 <= my_rom(2548); 
 data3 <= my_rom(3903); 
 data4 <= my_rom(5258); 
 data5 <= my_rom(6613); 
 data6 <= my_rom(7968); 
 data7 <= my_rom(9323); 
 data8 <= my_rom(10678); 
 data9 <= my_rom(12033); 
 data10 <= my_rom(13388);
when "10010101010" => 
 data1 <= my_rom(1194); 
 data2 <= my_rom(2549); 
 data3 <= my_rom(3904); 
 data4 <= my_rom(5259); 
 data5 <= my_rom(6614); 
 data6 <= my_rom(7969); 
 data7 <= my_rom(9324); 
 data8 <= my_rom(10679); 
 data9 <= my_rom(12034); 
 data10 <= my_rom(13389);
when "10010101011" => 
 data1 <= my_rom(1195); 
 data2 <= my_rom(2550); 
 data3 <= my_rom(3905); 
 data4 <= my_rom(5260); 
 data5 <= my_rom(6615); 
 data6 <= my_rom(7970); 
 data7 <= my_rom(9325); 
 data8 <= my_rom(10680); 
 data9 <= my_rom(12035); 
 data10 <= my_rom(13390);
when "10010101100" => 
 data1 <= my_rom(1196); 
 data2 <= my_rom(2551); 
 data3 <= my_rom(3906); 
 data4 <= my_rom(5261); 
 data5 <= my_rom(6616); 
 data6 <= my_rom(7971); 
 data7 <= my_rom(9326); 
 data8 <= my_rom(10681); 
 data9 <= my_rom(12036); 
 data10 <= my_rom(13391);
when "10010101101" => 
 data1 <= my_rom(1197); 
 data2 <= my_rom(2552); 
 data3 <= my_rom(3907); 
 data4 <= my_rom(5262); 
 data5 <= my_rom(6617); 
 data6 <= my_rom(7972); 
 data7 <= my_rom(9327); 
 data8 <= my_rom(10682); 
 data9 <= my_rom(12037); 
 data10 <= my_rom(13392);
when "10010101110" => 
 data1 <= my_rom(1198); 
 data2 <= my_rom(2553); 
 data3 <= my_rom(3908); 
 data4 <= my_rom(5263); 
 data5 <= my_rom(6618); 
 data6 <= my_rom(7973); 
 data7 <= my_rom(9328); 
 data8 <= my_rom(10683); 
 data9 <= my_rom(12038); 
 data10 <= my_rom(13393);
when "10010101111" => 
 data1 <= my_rom(1199); 
 data2 <= my_rom(2554); 
 data3 <= my_rom(3909); 
 data4 <= my_rom(5264); 
 data5 <= my_rom(6619); 
 data6 <= my_rom(7974); 
 data7 <= my_rom(9329); 
 data8 <= my_rom(10684); 
 data9 <= my_rom(12039); 
 data10 <= my_rom(13394);
when "10010110000" => 
 data1 <= my_rom(1200); 
 data2 <= my_rom(2555); 
 data3 <= my_rom(3910); 
 data4 <= my_rom(5265); 
 data5 <= my_rom(6620); 
 data6 <= my_rom(7975); 
 data7 <= my_rom(9330); 
 data8 <= my_rom(10685); 
 data9 <= my_rom(12040); 
 data10 <= my_rom(13395);
when "10010110001" => 
 data1 <= my_rom(1201); 
 data2 <= my_rom(2556); 
 data3 <= my_rom(3911); 
 data4 <= my_rom(5266); 
 data5 <= my_rom(6621); 
 data6 <= my_rom(7976); 
 data7 <= my_rom(9331); 
 data8 <= my_rom(10686); 
 data9 <= my_rom(12041); 
 data10 <= my_rom(13396);
when "10010110010" => 
 data1 <= my_rom(1202); 
 data2 <= my_rom(2557); 
 data3 <= my_rom(3912); 
 data4 <= my_rom(5267); 
 data5 <= my_rom(6622); 
 data6 <= my_rom(7977); 
 data7 <= my_rom(9332); 
 data8 <= my_rom(10687); 
 data9 <= my_rom(12042); 
 data10 <= my_rom(13397);
when "10010110011" => 
 data1 <= my_rom(1203); 
 data2 <= my_rom(2558); 
 data3 <= my_rom(3913); 
 data4 <= my_rom(5268); 
 data5 <= my_rom(6623); 
 data6 <= my_rom(7978); 
 data7 <= my_rom(9333); 
 data8 <= my_rom(10688); 
 data9 <= my_rom(12043); 
 data10 <= my_rom(13398);
when "10010110100" => 
 data1 <= my_rom(1204); 
 data2 <= my_rom(2559); 
 data3 <= my_rom(3914); 
 data4 <= my_rom(5269); 
 data5 <= my_rom(6624); 
 data6 <= my_rom(7979); 
 data7 <= my_rom(9334); 
 data8 <= my_rom(10689); 
 data9 <= my_rom(12044); 
 data10 <= my_rom(13399);
when "10010110101" => 
 data1 <= my_rom(1205); 
 data2 <= my_rom(2560); 
 data3 <= my_rom(3915); 
 data4 <= my_rom(5270); 
 data5 <= my_rom(6625); 
 data6 <= my_rom(7980); 
 data7 <= my_rom(9335); 
 data8 <= my_rom(10690); 
 data9 <= my_rom(12045); 
 data10 <= my_rom(13400);
when "10010110110" => 
 data1 <= my_rom(1206); 
 data2 <= my_rom(2561); 
 data3 <= my_rom(3916); 
 data4 <= my_rom(5271); 
 data5 <= my_rom(6626); 
 data6 <= my_rom(7981); 
 data7 <= my_rom(9336); 
 data8 <= my_rom(10691); 
 data9 <= my_rom(12046); 
 data10 <= my_rom(13401);
when "10010110111" => 
 data1 <= my_rom(1207); 
 data2 <= my_rom(2562); 
 data3 <= my_rom(3917); 
 data4 <= my_rom(5272); 
 data5 <= my_rom(6627); 
 data6 <= my_rom(7982); 
 data7 <= my_rom(9337); 
 data8 <= my_rom(10692); 
 data9 <= my_rom(12047); 
 data10 <= my_rom(13402);
when "10010111000" => 
 data1 <= my_rom(1208); 
 data2 <= my_rom(2563); 
 data3 <= my_rom(3918); 
 data4 <= my_rom(5273); 
 data5 <= my_rom(6628); 
 data6 <= my_rom(7983); 
 data7 <= my_rom(9338); 
 data8 <= my_rom(10693); 
 data9 <= my_rom(12048); 
 data10 <= my_rom(13403);
when "10010111001" => 
 data1 <= my_rom(1209); 
 data2 <= my_rom(2564); 
 data3 <= my_rom(3919); 
 data4 <= my_rom(5274); 
 data5 <= my_rom(6629); 
 data6 <= my_rom(7984); 
 data7 <= my_rom(9339); 
 data8 <= my_rom(10694); 
 data9 <= my_rom(12049); 
 data10 <= my_rom(13404);
when "10010111010" => 
 data1 <= my_rom(1210); 
 data2 <= my_rom(2565); 
 data3 <= my_rom(3920); 
 data4 <= my_rom(5275); 
 data5 <= my_rom(6630); 
 data6 <= my_rom(7985); 
 data7 <= my_rom(9340); 
 data8 <= my_rom(10695); 
 data9 <= my_rom(12050); 
 data10 <= my_rom(13405);
when "10010111011" => 
 data1 <= my_rom(1211); 
 data2 <= my_rom(2566); 
 data3 <= my_rom(3921); 
 data4 <= my_rom(5276); 
 data5 <= my_rom(6631); 
 data6 <= my_rom(7986); 
 data7 <= my_rom(9341); 
 data8 <= my_rom(10696); 
 data9 <= my_rom(12051); 
 data10 <= my_rom(13406);
when "10010111100" => 
 data1 <= my_rom(1212); 
 data2 <= my_rom(2567); 
 data3 <= my_rom(3922); 
 data4 <= my_rom(5277); 
 data5 <= my_rom(6632); 
 data6 <= my_rom(7987); 
 data7 <= my_rom(9342); 
 data8 <= my_rom(10697); 
 data9 <= my_rom(12052); 
 data10 <= my_rom(13407);
when "10010111101" => 
 data1 <= my_rom(1213); 
 data2 <= my_rom(2568); 
 data3 <= my_rom(3923); 
 data4 <= my_rom(5278); 
 data5 <= my_rom(6633); 
 data6 <= my_rom(7988); 
 data7 <= my_rom(9343); 
 data8 <= my_rom(10698); 
 data9 <= my_rom(12053); 
 data10 <= my_rom(13408);
when "10010111110" => 
 data1 <= my_rom(1214); 
 data2 <= my_rom(2569); 
 data3 <= my_rom(3924); 
 data4 <= my_rom(5279); 
 data5 <= my_rom(6634); 
 data6 <= my_rom(7989); 
 data7 <= my_rom(9344); 
 data8 <= my_rom(10699); 
 data9 <= my_rom(12054); 
 data10 <= my_rom(13409);
when "10010111111" => 
 data1 <= my_rom(1215); 
 data2 <= my_rom(2570); 
 data3 <= my_rom(3925); 
 data4 <= my_rom(5280); 
 data5 <= my_rom(6635); 
 data6 <= my_rom(7990); 
 data7 <= my_rom(9345); 
 data8 <= my_rom(10700); 
 data9 <= my_rom(12055); 
 data10 <= my_rom(13410);
when "10011000000" => 
 data1 <= my_rom(1216); 
 data2 <= my_rom(2571); 
 data3 <= my_rom(3926); 
 data4 <= my_rom(5281); 
 data5 <= my_rom(6636); 
 data6 <= my_rom(7991); 
 data7 <= my_rom(9346); 
 data8 <= my_rom(10701); 
 data9 <= my_rom(12056); 
 data10 <= my_rom(13411);
when "10011000001" => 
 data1 <= my_rom(1217); 
 data2 <= my_rom(2572); 
 data3 <= my_rom(3927); 
 data4 <= my_rom(5282); 
 data5 <= my_rom(6637); 
 data6 <= my_rom(7992); 
 data7 <= my_rom(9347); 
 data8 <= my_rom(10702); 
 data9 <= my_rom(12057); 
 data10 <= my_rom(13412);
when "10011000010" => 
 data1 <= my_rom(1218); 
 data2 <= my_rom(2573); 
 data3 <= my_rom(3928); 
 data4 <= my_rom(5283); 
 data5 <= my_rom(6638); 
 data6 <= my_rom(7993); 
 data7 <= my_rom(9348); 
 data8 <= my_rom(10703); 
 data9 <= my_rom(12058); 
 data10 <= my_rom(13413);
when "10011000011" => 
 data1 <= my_rom(1219); 
 data2 <= my_rom(2574); 
 data3 <= my_rom(3929); 
 data4 <= my_rom(5284); 
 data5 <= my_rom(6639); 
 data6 <= my_rom(7994); 
 data7 <= my_rom(9349); 
 data8 <= my_rom(10704); 
 data9 <= my_rom(12059); 
 data10 <= my_rom(13414);
when "10011000100" => 
 data1 <= my_rom(1220); 
 data2 <= my_rom(2575); 
 data3 <= my_rom(3930); 
 data4 <= my_rom(5285); 
 data5 <= my_rom(6640); 
 data6 <= my_rom(7995); 
 data7 <= my_rom(9350); 
 data8 <= my_rom(10705); 
 data9 <= my_rom(12060); 
 data10 <= my_rom(13415);
when "10011000101" => 
 data1 <= my_rom(1221); 
 data2 <= my_rom(2576); 
 data3 <= my_rom(3931); 
 data4 <= my_rom(5286); 
 data5 <= my_rom(6641); 
 data6 <= my_rom(7996); 
 data7 <= my_rom(9351); 
 data8 <= my_rom(10706); 
 data9 <= my_rom(12061); 
 data10 <= my_rom(13416);
when "10011000110" => 
 data1 <= my_rom(1222); 
 data2 <= my_rom(2577); 
 data3 <= my_rom(3932); 
 data4 <= my_rom(5287); 
 data5 <= my_rom(6642); 
 data6 <= my_rom(7997); 
 data7 <= my_rom(9352); 
 data8 <= my_rom(10707); 
 data9 <= my_rom(12062); 
 data10 <= my_rom(13417);
when "10011000111" => 
 data1 <= my_rom(1223); 
 data2 <= my_rom(2578); 
 data3 <= my_rom(3933); 
 data4 <= my_rom(5288); 
 data5 <= my_rom(6643); 
 data6 <= my_rom(7998); 
 data7 <= my_rom(9353); 
 data8 <= my_rom(10708); 
 data9 <= my_rom(12063); 
 data10 <= my_rom(13418);
when "10011001000" => 
 data1 <= my_rom(1224); 
 data2 <= my_rom(2579); 
 data3 <= my_rom(3934); 
 data4 <= my_rom(5289); 
 data5 <= my_rom(6644); 
 data6 <= my_rom(7999); 
 data7 <= my_rom(9354); 
 data8 <= my_rom(10709); 
 data9 <= my_rom(12064); 
 data10 <= my_rom(13419);
when "10011001001" => 
 data1 <= my_rom(1225); 
 data2 <= my_rom(2580); 
 data3 <= my_rom(3935); 
 data4 <= my_rom(5290); 
 data5 <= my_rom(6645); 
 data6 <= my_rom(8000); 
 data7 <= my_rom(9355); 
 data8 <= my_rom(10710); 
 data9 <= my_rom(12065); 
 data10 <= my_rom(13420);
when "10011001010" => 
 data1 <= my_rom(1226); 
 data2 <= my_rom(2581); 
 data3 <= my_rom(3936); 
 data4 <= my_rom(5291); 
 data5 <= my_rom(6646); 
 data6 <= my_rom(8001); 
 data7 <= my_rom(9356); 
 data8 <= my_rom(10711); 
 data9 <= my_rom(12066); 
 data10 <= my_rom(13421);
when "10011001011" => 
 data1 <= my_rom(1227); 
 data2 <= my_rom(2582); 
 data3 <= my_rom(3937); 
 data4 <= my_rom(5292); 
 data5 <= my_rom(6647); 
 data6 <= my_rom(8002); 
 data7 <= my_rom(9357); 
 data8 <= my_rom(10712); 
 data9 <= my_rom(12067); 
 data10 <= my_rom(13422);
when "10011001100" => 
 data1 <= my_rom(1228); 
 data2 <= my_rom(2583); 
 data3 <= my_rom(3938); 
 data4 <= my_rom(5293); 
 data5 <= my_rom(6648); 
 data6 <= my_rom(8003); 
 data7 <= my_rom(9358); 
 data8 <= my_rom(10713); 
 data9 <= my_rom(12068); 
 data10 <= my_rom(13423);
when "10011001101" => 
 data1 <= my_rom(1229); 
 data2 <= my_rom(2584); 
 data3 <= my_rom(3939); 
 data4 <= my_rom(5294); 
 data5 <= my_rom(6649); 
 data6 <= my_rom(8004); 
 data7 <= my_rom(9359); 
 data8 <= my_rom(10714); 
 data9 <= my_rom(12069); 
 data10 <= my_rom(13424);
when "10011001110" => 
 data1 <= my_rom(1230); 
 data2 <= my_rom(2585); 
 data3 <= my_rom(3940); 
 data4 <= my_rom(5295); 
 data5 <= my_rom(6650); 
 data6 <= my_rom(8005); 
 data7 <= my_rom(9360); 
 data8 <= my_rom(10715); 
 data9 <= my_rom(12070); 
 data10 <= my_rom(13425);
when "10011001111" => 
 data1 <= my_rom(1231); 
 data2 <= my_rom(2586); 
 data3 <= my_rom(3941); 
 data4 <= my_rom(5296); 
 data5 <= my_rom(6651); 
 data6 <= my_rom(8006); 
 data7 <= my_rom(9361); 
 data8 <= my_rom(10716); 
 data9 <= my_rom(12071); 
 data10 <= my_rom(13426);
when "10011010000" => 
 data1 <= my_rom(1232); 
 data2 <= my_rom(2587); 
 data3 <= my_rom(3942); 
 data4 <= my_rom(5297); 
 data5 <= my_rom(6652); 
 data6 <= my_rom(8007); 
 data7 <= my_rom(9362); 
 data8 <= my_rom(10717); 
 data9 <= my_rom(12072); 
 data10 <= my_rom(13427);
when "10011010001" => 
 data1 <= my_rom(1233); 
 data2 <= my_rom(2588); 
 data3 <= my_rom(3943); 
 data4 <= my_rom(5298); 
 data5 <= my_rom(6653); 
 data6 <= my_rom(8008); 
 data7 <= my_rom(9363); 
 data8 <= my_rom(10718); 
 data9 <= my_rom(12073); 
 data10 <= my_rom(13428);
when "10011010010" => 
 data1 <= my_rom(1234); 
 data2 <= my_rom(2589); 
 data3 <= my_rom(3944); 
 data4 <= my_rom(5299); 
 data5 <= my_rom(6654); 
 data6 <= my_rom(8009); 
 data7 <= my_rom(9364); 
 data8 <= my_rom(10719); 
 data9 <= my_rom(12074); 
 data10 <= my_rom(13429);
when "10011010011" => 
 data1 <= my_rom(1235); 
 data2 <= my_rom(2590); 
 data3 <= my_rom(3945); 
 data4 <= my_rom(5300); 
 data5 <= my_rom(6655); 
 data6 <= my_rom(8010); 
 data7 <= my_rom(9365); 
 data8 <= my_rom(10720); 
 data9 <= my_rom(12075); 
 data10 <= my_rom(13430);
when "10011010100" => 
 data1 <= my_rom(1236); 
 data2 <= my_rom(2591); 
 data3 <= my_rom(3946); 
 data4 <= my_rom(5301); 
 data5 <= my_rom(6656); 
 data6 <= my_rom(8011); 
 data7 <= my_rom(9366); 
 data8 <= my_rom(10721); 
 data9 <= my_rom(12076); 
 data10 <= my_rom(13431);
when "10011010101" => 
 data1 <= my_rom(1237); 
 data2 <= my_rom(2592); 
 data3 <= my_rom(3947); 
 data4 <= my_rom(5302); 
 data5 <= my_rom(6657); 
 data6 <= my_rom(8012); 
 data7 <= my_rom(9367); 
 data8 <= my_rom(10722); 
 data9 <= my_rom(12077); 
 data10 <= my_rom(13432);
when "10011010110" => 
 data1 <= my_rom(1238); 
 data2 <= my_rom(2593); 
 data3 <= my_rom(3948); 
 data4 <= my_rom(5303); 
 data5 <= my_rom(6658); 
 data6 <= my_rom(8013); 
 data7 <= my_rom(9368); 
 data8 <= my_rom(10723); 
 data9 <= my_rom(12078); 
 data10 <= my_rom(13433);
when "10011010111" => 
 data1 <= my_rom(1239); 
 data2 <= my_rom(2594); 
 data3 <= my_rom(3949); 
 data4 <= my_rom(5304); 
 data5 <= my_rom(6659); 
 data6 <= my_rom(8014); 
 data7 <= my_rom(9369); 
 data8 <= my_rom(10724); 
 data9 <= my_rom(12079); 
 data10 <= my_rom(13434);
when "10011011000" => 
 data1 <= my_rom(1240); 
 data2 <= my_rom(2595); 
 data3 <= my_rom(3950); 
 data4 <= my_rom(5305); 
 data5 <= my_rom(6660); 
 data6 <= my_rom(8015); 
 data7 <= my_rom(9370); 
 data8 <= my_rom(10725); 
 data9 <= my_rom(12080); 
 data10 <= my_rom(13435);
when "10011011001" => 
 data1 <= my_rom(1241); 
 data2 <= my_rom(2596); 
 data3 <= my_rom(3951); 
 data4 <= my_rom(5306); 
 data5 <= my_rom(6661); 
 data6 <= my_rom(8016); 
 data7 <= my_rom(9371); 
 data8 <= my_rom(10726); 
 data9 <= my_rom(12081); 
 data10 <= my_rom(13436);
when "10011011010" => 
 data1 <= my_rom(1242); 
 data2 <= my_rom(2597); 
 data3 <= my_rom(3952); 
 data4 <= my_rom(5307); 
 data5 <= my_rom(6662); 
 data6 <= my_rom(8017); 
 data7 <= my_rom(9372); 
 data8 <= my_rom(10727); 
 data9 <= my_rom(12082); 
 data10 <= my_rom(13437);
when "10011011011" => 
 data1 <= my_rom(1243); 
 data2 <= my_rom(2598); 
 data3 <= my_rom(3953); 
 data4 <= my_rom(5308); 
 data5 <= my_rom(6663); 
 data6 <= my_rom(8018); 
 data7 <= my_rom(9373); 
 data8 <= my_rom(10728); 
 data9 <= my_rom(12083); 
 data10 <= my_rom(13438);
when "10011011100" => 
 data1 <= my_rom(1244); 
 data2 <= my_rom(2599); 
 data3 <= my_rom(3954); 
 data4 <= my_rom(5309); 
 data5 <= my_rom(6664); 
 data6 <= my_rom(8019); 
 data7 <= my_rom(9374); 
 data8 <= my_rom(10729); 
 data9 <= my_rom(12084); 
 data10 <= my_rom(13439);
when "10011011101" => 
 data1 <= my_rom(1245); 
 data2 <= my_rom(2600); 
 data3 <= my_rom(3955); 
 data4 <= my_rom(5310); 
 data5 <= my_rom(6665); 
 data6 <= my_rom(8020); 
 data7 <= my_rom(9375); 
 data8 <= my_rom(10730); 
 data9 <= my_rom(12085); 
 data10 <= my_rom(13440);
when "10011011110" => 
 data1 <= my_rom(1246); 
 data2 <= my_rom(2601); 
 data3 <= my_rom(3956); 
 data4 <= my_rom(5311); 
 data5 <= my_rom(6666); 
 data6 <= my_rom(8021); 
 data7 <= my_rom(9376); 
 data8 <= my_rom(10731); 
 data9 <= my_rom(12086); 
 data10 <= my_rom(13441);
when "10011011111" => 
 data1 <= my_rom(1247); 
 data2 <= my_rom(2602); 
 data3 <= my_rom(3957); 
 data4 <= my_rom(5312); 
 data5 <= my_rom(6667); 
 data6 <= my_rom(8022); 
 data7 <= my_rom(9377); 
 data8 <= my_rom(10732); 
 data9 <= my_rom(12087); 
 data10 <= my_rom(13442);
when "10011100000" => 
 data1 <= my_rom(1248); 
 data2 <= my_rom(2603); 
 data3 <= my_rom(3958); 
 data4 <= my_rom(5313); 
 data5 <= my_rom(6668); 
 data6 <= my_rom(8023); 
 data7 <= my_rom(9378); 
 data8 <= my_rom(10733); 
 data9 <= my_rom(12088); 
 data10 <= my_rom(13443);
when "10011100001" => 
 data1 <= my_rom(1249); 
 data2 <= my_rom(2604); 
 data3 <= my_rom(3959); 
 data4 <= my_rom(5314); 
 data5 <= my_rom(6669); 
 data6 <= my_rom(8024); 
 data7 <= my_rom(9379); 
 data8 <= my_rom(10734); 
 data9 <= my_rom(12089); 
 data10 <= my_rom(13444);
when "10011100010" => 
 data1 <= my_rom(1250); 
 data2 <= my_rom(2605); 
 data3 <= my_rom(3960); 
 data4 <= my_rom(5315); 
 data5 <= my_rom(6670); 
 data6 <= my_rom(8025); 
 data7 <= my_rom(9380); 
 data8 <= my_rom(10735); 
 data9 <= my_rom(12090); 
 data10 <= my_rom(13445);
when "10011100011" => 
 data1 <= my_rom(1251); 
 data2 <= my_rom(2606); 
 data3 <= my_rom(3961); 
 data4 <= my_rom(5316); 
 data5 <= my_rom(6671); 
 data6 <= my_rom(8026); 
 data7 <= my_rom(9381); 
 data8 <= my_rom(10736); 
 data9 <= my_rom(12091); 
 data10 <= my_rom(13446);
when "10011100100" => 
 data1 <= my_rom(1252); 
 data2 <= my_rom(2607); 
 data3 <= my_rom(3962); 
 data4 <= my_rom(5317); 
 data5 <= my_rom(6672); 
 data6 <= my_rom(8027); 
 data7 <= my_rom(9382); 
 data8 <= my_rom(10737); 
 data9 <= my_rom(12092); 
 data10 <= my_rom(13447);
when "10011100101" => 
 data1 <= my_rom(1253); 
 data2 <= my_rom(2608); 
 data3 <= my_rom(3963); 
 data4 <= my_rom(5318); 
 data5 <= my_rom(6673); 
 data6 <= my_rom(8028); 
 data7 <= my_rom(9383); 
 data8 <= my_rom(10738); 
 data9 <= my_rom(12093); 
 data10 <= my_rom(13448);
when "10011100110" => 
 data1 <= my_rom(1254); 
 data2 <= my_rom(2609); 
 data3 <= my_rom(3964); 
 data4 <= my_rom(5319); 
 data5 <= my_rom(6674); 
 data6 <= my_rom(8029); 
 data7 <= my_rom(9384); 
 data8 <= my_rom(10739); 
 data9 <= my_rom(12094); 
 data10 <= my_rom(13449);
when "10011100111" => 
 data1 <= my_rom(1255); 
 data2 <= my_rom(2610); 
 data3 <= my_rom(3965); 
 data4 <= my_rom(5320); 
 data5 <= my_rom(6675); 
 data6 <= my_rom(8030); 
 data7 <= my_rom(9385); 
 data8 <= my_rom(10740); 
 data9 <= my_rom(12095); 
 data10 <= my_rom(13450);
when "10011101000" => 
 data1 <= my_rom(1256); 
 data2 <= my_rom(2611); 
 data3 <= my_rom(3966); 
 data4 <= my_rom(5321); 
 data5 <= my_rom(6676); 
 data6 <= my_rom(8031); 
 data7 <= my_rom(9386); 
 data8 <= my_rom(10741); 
 data9 <= my_rom(12096); 
 data10 <= my_rom(13451);
when "10011101001" => 
 data1 <= my_rom(1257); 
 data2 <= my_rom(2612); 
 data3 <= my_rom(3967); 
 data4 <= my_rom(5322); 
 data5 <= my_rom(6677); 
 data6 <= my_rom(8032); 
 data7 <= my_rom(9387); 
 data8 <= my_rom(10742); 
 data9 <= my_rom(12097); 
 data10 <= my_rom(13452);
when "10011101010" => 
 data1 <= my_rom(1258); 
 data2 <= my_rom(2613); 
 data3 <= my_rom(3968); 
 data4 <= my_rom(5323); 
 data5 <= my_rom(6678); 
 data6 <= my_rom(8033); 
 data7 <= my_rom(9388); 
 data8 <= my_rom(10743); 
 data9 <= my_rom(12098); 
 data10 <= my_rom(13453);
when "10011101011" => 
 data1 <= my_rom(1259); 
 data2 <= my_rom(2614); 
 data3 <= my_rom(3969); 
 data4 <= my_rom(5324); 
 data5 <= my_rom(6679); 
 data6 <= my_rom(8034); 
 data7 <= my_rom(9389); 
 data8 <= my_rom(10744); 
 data9 <= my_rom(12099); 
 data10 <= my_rom(13454);
when "10011101100" => 
 data1 <= my_rom(1260); 
 data2 <= my_rom(2615); 
 data3 <= my_rom(3970); 
 data4 <= my_rom(5325); 
 data5 <= my_rom(6680); 
 data6 <= my_rom(8035); 
 data7 <= my_rom(9390); 
 data8 <= my_rom(10745); 
 data9 <= my_rom(12100); 
 data10 <= my_rom(13455);
when "10011101101" => 
 data1 <= my_rom(1261); 
 data2 <= my_rom(2616); 
 data3 <= my_rom(3971); 
 data4 <= my_rom(5326); 
 data5 <= my_rom(6681); 
 data6 <= my_rom(8036); 
 data7 <= my_rom(9391); 
 data8 <= my_rom(10746); 
 data9 <= my_rom(12101); 
 data10 <= my_rom(13456);
when "10011101110" => 
 data1 <= my_rom(1262); 
 data2 <= my_rom(2617); 
 data3 <= my_rom(3972); 
 data4 <= my_rom(5327); 
 data5 <= my_rom(6682); 
 data6 <= my_rom(8037); 
 data7 <= my_rom(9392); 
 data8 <= my_rom(10747); 
 data9 <= my_rom(12102); 
 data10 <= my_rom(13457);
when "10011101111" => 
 data1 <= my_rom(1263); 
 data2 <= my_rom(2618); 
 data3 <= my_rom(3973); 
 data4 <= my_rom(5328); 
 data5 <= my_rom(6683); 
 data6 <= my_rom(8038); 
 data7 <= my_rom(9393); 
 data8 <= my_rom(10748); 
 data9 <= my_rom(12103); 
 data10 <= my_rom(13458);
when "10011110000" => 
 data1 <= my_rom(1264); 
 data2 <= my_rom(2619); 
 data3 <= my_rom(3974); 
 data4 <= my_rom(5329); 
 data5 <= my_rom(6684); 
 data6 <= my_rom(8039); 
 data7 <= my_rom(9394); 
 data8 <= my_rom(10749); 
 data9 <= my_rom(12104); 
 data10 <= my_rom(13459);
when "10011110001" => 
 data1 <= my_rom(1265); 
 data2 <= my_rom(2620); 
 data3 <= my_rom(3975); 
 data4 <= my_rom(5330); 
 data5 <= my_rom(6685); 
 data6 <= my_rom(8040); 
 data7 <= my_rom(9395); 
 data8 <= my_rom(10750); 
 data9 <= my_rom(12105); 
 data10 <= my_rom(13460);
when "10011110010" => 
 data1 <= my_rom(1266); 
 data2 <= my_rom(2621); 
 data3 <= my_rom(3976); 
 data4 <= my_rom(5331); 
 data5 <= my_rom(6686); 
 data6 <= my_rom(8041); 
 data7 <= my_rom(9396); 
 data8 <= my_rom(10751); 
 data9 <= my_rom(12106); 
 data10 <= my_rom(13461);
when "10011110011" => 
 data1 <= my_rom(1267); 
 data2 <= my_rom(2622); 
 data3 <= my_rom(3977); 
 data4 <= my_rom(5332); 
 data5 <= my_rom(6687); 
 data6 <= my_rom(8042); 
 data7 <= my_rom(9397); 
 data8 <= my_rom(10752); 
 data9 <= my_rom(12107); 
 data10 <= my_rom(13462);
when "10011110100" => 
 data1 <= my_rom(1268); 
 data2 <= my_rom(2623); 
 data3 <= my_rom(3978); 
 data4 <= my_rom(5333); 
 data5 <= my_rom(6688); 
 data6 <= my_rom(8043); 
 data7 <= my_rom(9398); 
 data8 <= my_rom(10753); 
 data9 <= my_rom(12108); 
 data10 <= my_rom(13463);
when "10011110101" => 
 data1 <= my_rom(1269); 
 data2 <= my_rom(2624); 
 data3 <= my_rom(3979); 
 data4 <= my_rom(5334); 
 data5 <= my_rom(6689); 
 data6 <= my_rom(8044); 
 data7 <= my_rom(9399); 
 data8 <= my_rom(10754); 
 data9 <= my_rom(12109); 
 data10 <= my_rom(13464);
when "10011110110" => 
 data1 <= my_rom(1270); 
 data2 <= my_rom(2625); 
 data3 <= my_rom(3980); 
 data4 <= my_rom(5335); 
 data5 <= my_rom(6690); 
 data6 <= my_rom(8045); 
 data7 <= my_rom(9400); 
 data8 <= my_rom(10755); 
 data9 <= my_rom(12110); 
 data10 <= my_rom(13465);
when "10011110111" => 
 data1 <= my_rom(1271); 
 data2 <= my_rom(2626); 
 data3 <= my_rom(3981); 
 data4 <= my_rom(5336); 
 data5 <= my_rom(6691); 
 data6 <= my_rom(8046); 
 data7 <= my_rom(9401); 
 data8 <= my_rom(10756); 
 data9 <= my_rom(12111); 
 data10 <= my_rom(13466);
when "10011111000" => 
 data1 <= my_rom(1272); 
 data2 <= my_rom(2627); 
 data3 <= my_rom(3982); 
 data4 <= my_rom(5337); 
 data5 <= my_rom(6692); 
 data6 <= my_rom(8047); 
 data7 <= my_rom(9402); 
 data8 <= my_rom(10757); 
 data9 <= my_rom(12112); 
 data10 <= my_rom(13467);
when "10011111001" => 
 data1 <= my_rom(1273); 
 data2 <= my_rom(2628); 
 data3 <= my_rom(3983); 
 data4 <= my_rom(5338); 
 data5 <= my_rom(6693); 
 data6 <= my_rom(8048); 
 data7 <= my_rom(9403); 
 data8 <= my_rom(10758); 
 data9 <= my_rom(12113); 
 data10 <= my_rom(13468);
when "10011111010" => 
 data1 <= my_rom(1274); 
 data2 <= my_rom(2629); 
 data3 <= my_rom(3984); 
 data4 <= my_rom(5339); 
 data5 <= my_rom(6694); 
 data6 <= my_rom(8049); 
 data7 <= my_rom(9404); 
 data8 <= my_rom(10759); 
 data9 <= my_rom(12114); 
 data10 <= my_rom(13469);
when "10011111011" => 
 data1 <= my_rom(1275); 
 data2 <= my_rom(2630); 
 data3 <= my_rom(3985); 
 data4 <= my_rom(5340); 
 data5 <= my_rom(6695); 
 data6 <= my_rom(8050); 
 data7 <= my_rom(9405); 
 data8 <= my_rom(10760); 
 data9 <= my_rom(12115); 
 data10 <= my_rom(13470);
when "10011111100" => 
 data1 <= my_rom(1276); 
 data2 <= my_rom(2631); 
 data3 <= my_rom(3986); 
 data4 <= my_rom(5341); 
 data5 <= my_rom(6696); 
 data6 <= my_rom(8051); 
 data7 <= my_rom(9406); 
 data8 <= my_rom(10761); 
 data9 <= my_rom(12116); 
 data10 <= my_rom(13471);
when "10011111101" => 
 data1 <= my_rom(1277); 
 data2 <= my_rom(2632); 
 data3 <= my_rom(3987); 
 data4 <= my_rom(5342); 
 data5 <= my_rom(6697); 
 data6 <= my_rom(8052); 
 data7 <= my_rom(9407); 
 data8 <= my_rom(10762); 
 data9 <= my_rom(12117); 
 data10 <= my_rom(13472);
when "10011111110" => 
 data1 <= my_rom(1278); 
 data2 <= my_rom(2633); 
 data3 <= my_rom(3988); 
 data4 <= my_rom(5343); 
 data5 <= my_rom(6698); 
 data6 <= my_rom(8053); 
 data7 <= my_rom(9408); 
 data8 <= my_rom(10763); 
 data9 <= my_rom(12118); 
 data10 <= my_rom(13473);
when "10011111111" => 
 data1 <= my_rom(1279); 
 data2 <= my_rom(2634); 
 data3 <= my_rom(3989); 
 data4 <= my_rom(5344); 
 data5 <= my_rom(6699); 
 data6 <= my_rom(8054); 
 data7 <= my_rom(9409); 
 data8 <= my_rom(10764); 
 data9 <= my_rom(12119); 
 data10 <= my_rom(13474);
when "10100000000" => 
 data1 <= my_rom(1280); 
 data2 <= my_rom(2635); 
 data3 <= my_rom(3990); 
 data4 <= my_rom(5345); 
 data5 <= my_rom(6700); 
 data6 <= my_rom(8055); 
 data7 <= my_rom(9410); 
 data8 <= my_rom(10765); 
 data9 <= my_rom(12120); 
 data10 <= my_rom(13475);
when "10100000001" => 
 data1 <= my_rom(1281); 
 data2 <= my_rom(2636); 
 data3 <= my_rom(3991); 
 data4 <= my_rom(5346); 
 data5 <= my_rom(6701); 
 data6 <= my_rom(8056); 
 data7 <= my_rom(9411); 
 data8 <= my_rom(10766); 
 data9 <= my_rom(12121); 
 data10 <= my_rom(13476);
when "10100000010" => 
 data1 <= my_rom(1282); 
 data2 <= my_rom(2637); 
 data3 <= my_rom(3992); 
 data4 <= my_rom(5347); 
 data5 <= my_rom(6702); 
 data6 <= my_rom(8057); 
 data7 <= my_rom(9412); 
 data8 <= my_rom(10767); 
 data9 <= my_rom(12122); 
 data10 <= my_rom(13477);
when "10100000011" => 
 data1 <= my_rom(1283); 
 data2 <= my_rom(2638); 
 data3 <= my_rom(3993); 
 data4 <= my_rom(5348); 
 data5 <= my_rom(6703); 
 data6 <= my_rom(8058); 
 data7 <= my_rom(9413); 
 data8 <= my_rom(10768); 
 data9 <= my_rom(12123); 
 data10 <= my_rom(13478);
when "10100000100" => 
 data1 <= my_rom(1284); 
 data2 <= my_rom(2639); 
 data3 <= my_rom(3994); 
 data4 <= my_rom(5349); 
 data5 <= my_rom(6704); 
 data6 <= my_rom(8059); 
 data7 <= my_rom(9414); 
 data8 <= my_rom(10769); 
 data9 <= my_rom(12124); 
 data10 <= my_rom(13479);
when "10100000101" => 
 data1 <= my_rom(1285); 
 data2 <= my_rom(2640); 
 data3 <= my_rom(3995); 
 data4 <= my_rom(5350); 
 data5 <= my_rom(6705); 
 data6 <= my_rom(8060); 
 data7 <= my_rom(9415); 
 data8 <= my_rom(10770); 
 data9 <= my_rom(12125); 
 data10 <= my_rom(13480);
when "10100000110" => 
 data1 <= my_rom(1286); 
 data2 <= my_rom(2641); 
 data3 <= my_rom(3996); 
 data4 <= my_rom(5351); 
 data5 <= my_rom(6706); 
 data6 <= my_rom(8061); 
 data7 <= my_rom(9416); 
 data8 <= my_rom(10771); 
 data9 <= my_rom(12126); 
 data10 <= my_rom(13481);
when "10100000111" => 
 data1 <= my_rom(1287); 
 data2 <= my_rom(2642); 
 data3 <= my_rom(3997); 
 data4 <= my_rom(5352); 
 data5 <= my_rom(6707); 
 data6 <= my_rom(8062); 
 data7 <= my_rom(9417); 
 data8 <= my_rom(10772); 
 data9 <= my_rom(12127); 
 data10 <= my_rom(13482);
when "10100001000" => 
 data1 <= my_rom(1288); 
 data2 <= my_rom(2643); 
 data3 <= my_rom(3998); 
 data4 <= my_rom(5353); 
 data5 <= my_rom(6708); 
 data6 <= my_rom(8063); 
 data7 <= my_rom(9418); 
 data8 <= my_rom(10773); 
 data9 <= my_rom(12128); 
 data10 <= my_rom(13483);
when "10100001001" => 
 data1 <= my_rom(1289); 
 data2 <= my_rom(2644); 
 data3 <= my_rom(3999); 
 data4 <= my_rom(5354); 
 data5 <= my_rom(6709); 
 data6 <= my_rom(8064); 
 data7 <= my_rom(9419); 
 data8 <= my_rom(10774); 
 data9 <= my_rom(12129); 
 data10 <= my_rom(13484);
when "10100001010" => 
 data1 <= my_rom(1290); 
 data2 <= my_rom(2645); 
 data3 <= my_rom(4000); 
 data4 <= my_rom(5355); 
 data5 <= my_rom(6710); 
 data6 <= my_rom(8065); 
 data7 <= my_rom(9420); 
 data8 <= my_rom(10775); 
 data9 <= my_rom(12130); 
 data10 <= my_rom(13485);
when "10100001011" => 
 data1 <= my_rom(1291); 
 data2 <= my_rom(2646); 
 data3 <= my_rom(4001); 
 data4 <= my_rom(5356); 
 data5 <= my_rom(6711); 
 data6 <= my_rom(8066); 
 data7 <= my_rom(9421); 
 data8 <= my_rom(10776); 
 data9 <= my_rom(12131); 
 data10 <= my_rom(13486);
when "10100001100" => 
 data1 <= my_rom(1292); 
 data2 <= my_rom(2647); 
 data3 <= my_rom(4002); 
 data4 <= my_rom(5357); 
 data5 <= my_rom(6712); 
 data6 <= my_rom(8067); 
 data7 <= my_rom(9422); 
 data8 <= my_rom(10777); 
 data9 <= my_rom(12132); 
 data10 <= my_rom(13487);
when "10100001101" => 
 data1 <= my_rom(1293); 
 data2 <= my_rom(2648); 
 data3 <= my_rom(4003); 
 data4 <= my_rom(5358); 
 data5 <= my_rom(6713); 
 data6 <= my_rom(8068); 
 data7 <= my_rom(9423); 
 data8 <= my_rom(10778); 
 data9 <= my_rom(12133); 
 data10 <= my_rom(13488);
when "10100001110" => 
 data1 <= my_rom(1294); 
 data2 <= my_rom(2649); 
 data3 <= my_rom(4004); 
 data4 <= my_rom(5359); 
 data5 <= my_rom(6714); 
 data6 <= my_rom(8069); 
 data7 <= my_rom(9424); 
 data8 <= my_rom(10779); 
 data9 <= my_rom(12134); 
 data10 <= my_rom(13489);
when "10100001111" => 
 data1 <= my_rom(1295); 
 data2 <= my_rom(2650); 
 data3 <= my_rom(4005); 
 data4 <= my_rom(5360); 
 data5 <= my_rom(6715); 
 data6 <= my_rom(8070); 
 data7 <= my_rom(9425); 
 data8 <= my_rom(10780); 
 data9 <= my_rom(12135); 
 data10 <= my_rom(13490);
when "10100010000" => 
 data1 <= my_rom(1296); 
 data2 <= my_rom(2651); 
 data3 <= my_rom(4006); 
 data4 <= my_rom(5361); 
 data5 <= my_rom(6716); 
 data6 <= my_rom(8071); 
 data7 <= my_rom(9426); 
 data8 <= my_rom(10781); 
 data9 <= my_rom(12136); 
 data10 <= my_rom(13491);
when "10100010001" => 
 data1 <= my_rom(1297); 
 data2 <= my_rom(2652); 
 data3 <= my_rom(4007); 
 data4 <= my_rom(5362); 
 data5 <= my_rom(6717); 
 data6 <= my_rom(8072); 
 data7 <= my_rom(9427); 
 data8 <= my_rom(10782); 
 data9 <= my_rom(12137); 
 data10 <= my_rom(13492);
when "10100010010" => 
 data1 <= my_rom(1298); 
 data2 <= my_rom(2653); 
 data3 <= my_rom(4008); 
 data4 <= my_rom(5363); 
 data5 <= my_rom(6718); 
 data6 <= my_rom(8073); 
 data7 <= my_rom(9428); 
 data8 <= my_rom(10783); 
 data9 <= my_rom(12138); 
 data10 <= my_rom(13493);
when "10100010011" => 
 data1 <= my_rom(1299); 
 data2 <= my_rom(2654); 
 data3 <= my_rom(4009); 
 data4 <= my_rom(5364); 
 data5 <= my_rom(6719); 
 data6 <= my_rom(8074); 
 data7 <= my_rom(9429); 
 data8 <= my_rom(10784); 
 data9 <= my_rom(12139); 
 data10 <= my_rom(13494);
when "10100010100" => 
 data1 <= my_rom(1300); 
 data2 <= my_rom(2655); 
 data3 <= my_rom(4010); 
 data4 <= my_rom(5365); 
 data5 <= my_rom(6720); 
 data6 <= my_rom(8075); 
 data7 <= my_rom(9430); 
 data8 <= my_rom(10785); 
 data9 <= my_rom(12140); 
 data10 <= my_rom(13495);
when "10100010101" => 
 data1 <= my_rom(1301); 
 data2 <= my_rom(2656); 
 data3 <= my_rom(4011); 
 data4 <= my_rom(5366); 
 data5 <= my_rom(6721); 
 data6 <= my_rom(8076); 
 data7 <= my_rom(9431); 
 data8 <= my_rom(10786); 
 data9 <= my_rom(12141); 
 data10 <= my_rom(13496);
when "10100010110" => 
 data1 <= my_rom(1302); 
 data2 <= my_rom(2657); 
 data3 <= my_rom(4012); 
 data4 <= my_rom(5367); 
 data5 <= my_rom(6722); 
 data6 <= my_rom(8077); 
 data7 <= my_rom(9432); 
 data8 <= my_rom(10787); 
 data9 <= my_rom(12142); 
 data10 <= my_rom(13497);
when "10100010111" => 
 data1 <= my_rom(1303); 
 data2 <= my_rom(2658); 
 data3 <= my_rom(4013); 
 data4 <= my_rom(5368); 
 data5 <= my_rom(6723); 
 data6 <= my_rom(8078); 
 data7 <= my_rom(9433); 
 data8 <= my_rom(10788); 
 data9 <= my_rom(12143); 
 data10 <= my_rom(13498);
when "10100011000" => 
 data1 <= my_rom(1304); 
 data2 <= my_rom(2659); 
 data3 <= my_rom(4014); 
 data4 <= my_rom(5369); 
 data5 <= my_rom(6724); 
 data6 <= my_rom(8079); 
 data7 <= my_rom(9434); 
 data8 <= my_rom(10789); 
 data9 <= my_rom(12144); 
 data10 <= my_rom(13499);
when "10100011001" => 
 data1 <= my_rom(1305); 
 data2 <= my_rom(2660); 
 data3 <= my_rom(4015); 
 data4 <= my_rom(5370); 
 data5 <= my_rom(6725); 
 data6 <= my_rom(8080); 
 data7 <= my_rom(9435); 
 data8 <= my_rom(10790); 
 data9 <= my_rom(12145); 
 data10 <= my_rom(13500);
when "10100011010" => 
 data1 <= my_rom(1306); 
 data2 <= my_rom(2661); 
 data3 <= my_rom(4016); 
 data4 <= my_rom(5371); 
 data5 <= my_rom(6726); 
 data6 <= my_rom(8081); 
 data7 <= my_rom(9436); 
 data8 <= my_rom(10791); 
 data9 <= my_rom(12146); 
 data10 <= my_rom(13501);
when "10100011011" => 
 data1 <= my_rom(1307); 
 data2 <= my_rom(2662); 
 data3 <= my_rom(4017); 
 data4 <= my_rom(5372); 
 data5 <= my_rom(6727); 
 data6 <= my_rom(8082); 
 data7 <= my_rom(9437); 
 data8 <= my_rom(10792); 
 data9 <= my_rom(12147); 
 data10 <= my_rom(13502);
when "10100011100" => 
 data1 <= my_rom(1308); 
 data2 <= my_rom(2663); 
 data3 <= my_rom(4018); 
 data4 <= my_rom(5373); 
 data5 <= my_rom(6728); 
 data6 <= my_rom(8083); 
 data7 <= my_rom(9438); 
 data8 <= my_rom(10793); 
 data9 <= my_rom(12148); 
 data10 <= my_rom(13503);
when "10100011101" => 
 data1 <= my_rom(1309); 
 data2 <= my_rom(2664); 
 data3 <= my_rom(4019); 
 data4 <= my_rom(5374); 
 data5 <= my_rom(6729); 
 data6 <= my_rom(8084); 
 data7 <= my_rom(9439); 
 data8 <= my_rom(10794); 
 data9 <= my_rom(12149); 
 data10 <= my_rom(13504);
when "10100011110" => 
 data1 <= my_rom(1310); 
 data2 <= my_rom(2665); 
 data3 <= my_rom(4020); 
 data4 <= my_rom(5375); 
 data5 <= my_rom(6730); 
 data6 <= my_rom(8085); 
 data7 <= my_rom(9440); 
 data8 <= my_rom(10795); 
 data9 <= my_rom(12150); 
 data10 <= my_rom(13505);
when "10100011111" => 
 data1 <= my_rom(1311); 
 data2 <= my_rom(2666); 
 data3 <= my_rom(4021); 
 data4 <= my_rom(5376); 
 data5 <= my_rom(6731); 
 data6 <= my_rom(8086); 
 data7 <= my_rom(9441); 
 data8 <= my_rom(10796); 
 data9 <= my_rom(12151); 
 data10 <= my_rom(13506);
when "10100100000" => 
 data1 <= my_rom(1312); 
 data2 <= my_rom(2667); 
 data3 <= my_rom(4022); 
 data4 <= my_rom(5377); 
 data5 <= my_rom(6732); 
 data6 <= my_rom(8087); 
 data7 <= my_rom(9442); 
 data8 <= my_rom(10797); 
 data9 <= my_rom(12152); 
 data10 <= my_rom(13507);
when "10100100001" => 
 data1 <= my_rom(1313); 
 data2 <= my_rom(2668); 
 data3 <= my_rom(4023); 
 data4 <= my_rom(5378); 
 data5 <= my_rom(6733); 
 data6 <= my_rom(8088); 
 data7 <= my_rom(9443); 
 data8 <= my_rom(10798); 
 data9 <= my_rom(12153); 
 data10 <= my_rom(13508);
when "10100100010" => 
 data1 <= my_rom(1314); 
 data2 <= my_rom(2669); 
 data3 <= my_rom(4024); 
 data4 <= my_rom(5379); 
 data5 <= my_rom(6734); 
 data6 <= my_rom(8089); 
 data7 <= my_rom(9444); 
 data8 <= my_rom(10799); 
 data9 <= my_rom(12154); 
 data10 <= my_rom(13509);
when "10100100011" => 
 data1 <= my_rom(1315); 
 data2 <= my_rom(2670); 
 data3 <= my_rom(4025); 
 data4 <= my_rom(5380); 
 data5 <= my_rom(6735); 
 data6 <= my_rom(8090); 
 data7 <= my_rom(9445); 
 data8 <= my_rom(10800); 
 data9 <= my_rom(12155); 
 data10 <= my_rom(13510);
when "10100100100" => 
 data1 <= my_rom(1316); 
 data2 <= my_rom(2671); 
 data3 <= my_rom(4026); 
 data4 <= my_rom(5381); 
 data5 <= my_rom(6736); 
 data6 <= my_rom(8091); 
 data7 <= my_rom(9446); 
 data8 <= my_rom(10801); 
 data9 <= my_rom(12156); 
 data10 <= my_rom(13511);
when "10100100101" => 
 data1 <= my_rom(1317); 
 data2 <= my_rom(2672); 
 data3 <= my_rom(4027); 
 data4 <= my_rom(5382); 
 data5 <= my_rom(6737); 
 data6 <= my_rom(8092); 
 data7 <= my_rom(9447); 
 data8 <= my_rom(10802); 
 data9 <= my_rom(12157); 
 data10 <= my_rom(13512);
when "10100100110" => 
 data1 <= my_rom(1318); 
 data2 <= my_rom(2673); 
 data3 <= my_rom(4028); 
 data4 <= my_rom(5383); 
 data5 <= my_rom(6738); 
 data6 <= my_rom(8093); 
 data7 <= my_rom(9448); 
 data8 <= my_rom(10803); 
 data9 <= my_rom(12158); 
 data10 <= my_rom(13513);
when "10100100111" => 
 data1 <= my_rom(1319); 
 data2 <= my_rom(2674); 
 data3 <= my_rom(4029); 
 data4 <= my_rom(5384); 
 data5 <= my_rom(6739); 
 data6 <= my_rom(8094); 
 data7 <= my_rom(9449); 
 data8 <= my_rom(10804); 
 data9 <= my_rom(12159); 
 data10 <= my_rom(13514);
when "10100101000" => 
 data1 <= my_rom(1320); 
 data2 <= my_rom(2675); 
 data3 <= my_rom(4030); 
 data4 <= my_rom(5385); 
 data5 <= my_rom(6740); 
 data6 <= my_rom(8095); 
 data7 <= my_rom(9450); 
 data8 <= my_rom(10805); 
 data9 <= my_rom(12160); 
 data10 <= my_rom(13515);
when "10100101001" => 
 data1 <= my_rom(1321); 
 data2 <= my_rom(2676); 
 data3 <= my_rom(4031); 
 data4 <= my_rom(5386); 
 data5 <= my_rom(6741); 
 data6 <= my_rom(8096); 
 data7 <= my_rom(9451); 
 data8 <= my_rom(10806); 
 data9 <= my_rom(12161); 
 data10 <= my_rom(13516);
when "10100101010" => 
 data1 <= my_rom(1322); 
 data2 <= my_rom(2677); 
 data3 <= my_rom(4032); 
 data4 <= my_rom(5387); 
 data5 <= my_rom(6742); 
 data6 <= my_rom(8097); 
 data7 <= my_rom(9452); 
 data8 <= my_rom(10807); 
 data9 <= my_rom(12162); 
 data10 <= my_rom(13517);
when "10100101011" => 
 data1 <= my_rom(1323); 
 data2 <= my_rom(2678); 
 data3 <= my_rom(4033); 
 data4 <= my_rom(5388); 
 data5 <= my_rom(6743); 
 data6 <= my_rom(8098); 
 data7 <= my_rom(9453); 
 data8 <= my_rom(10808); 
 data9 <= my_rom(12163); 
 data10 <= my_rom(13518);
when "10100101100" => 
 data1 <= my_rom(1324); 
 data2 <= my_rom(2679); 
 data3 <= my_rom(4034); 
 data4 <= my_rom(5389); 
 data5 <= my_rom(6744); 
 data6 <= my_rom(8099); 
 data7 <= my_rom(9454); 
 data8 <= my_rom(10809); 
 data9 <= my_rom(12164); 
 data10 <= my_rom(13519);
when "10100101101" => 
 data1 <= my_rom(1325); 
 data2 <= my_rom(2680); 
 data3 <= my_rom(4035); 
 data4 <= my_rom(5390); 
 data5 <= my_rom(6745); 
 data6 <= my_rom(8100); 
 data7 <= my_rom(9455); 
 data8 <= my_rom(10810); 
 data9 <= my_rom(12165); 
 data10 <= my_rom(13520);
when "10100101110" => 
 data1 <= my_rom(1326); 
 data2 <= my_rom(2681); 
 data3 <= my_rom(4036); 
 data4 <= my_rom(5391); 
 data5 <= my_rom(6746); 
 data6 <= my_rom(8101); 
 data7 <= my_rom(9456); 
 data8 <= my_rom(10811); 
 data9 <= my_rom(12166); 
 data10 <= my_rom(13521);
when "10100101111" => 
 data1 <= my_rom(1327); 
 data2 <= my_rom(2682); 
 data3 <= my_rom(4037); 
 data4 <= my_rom(5392); 
 data5 <= my_rom(6747); 
 data6 <= my_rom(8102); 
 data7 <= my_rom(9457); 
 data8 <= my_rom(10812); 
 data9 <= my_rom(12167); 
 data10 <= my_rom(13522);
when "10100110000" => 
 data1 <= my_rom(1328); 
 data2 <= my_rom(2683); 
 data3 <= my_rom(4038); 
 data4 <= my_rom(5393); 
 data5 <= my_rom(6748); 
 data6 <= my_rom(8103); 
 data7 <= my_rom(9458); 
 data8 <= my_rom(10813); 
 data9 <= my_rom(12168); 
 data10 <= my_rom(13523);
when "10100110001" => 
 data1 <= my_rom(1329); 
 data2 <= my_rom(2684); 
 data3 <= my_rom(4039); 
 data4 <= my_rom(5394); 
 data5 <= my_rom(6749); 
 data6 <= my_rom(8104); 
 data7 <= my_rom(9459); 
 data8 <= my_rom(10814); 
 data9 <= my_rom(12169); 
 data10 <= my_rom(13524);
when "10100110010" => 
 data1 <= my_rom(1330); 
 data2 <= my_rom(2685); 
 data3 <= my_rom(4040); 
 data4 <= my_rom(5395); 
 data5 <= my_rom(6750); 
 data6 <= my_rom(8105); 
 data7 <= my_rom(9460); 
 data8 <= my_rom(10815); 
 data9 <= my_rom(12170); 
 data10 <= my_rom(13525);
when "10100110011" => 
 data1 <= my_rom(1331); 
 data2 <= my_rom(2686); 
 data3 <= my_rom(4041); 
 data4 <= my_rom(5396); 
 data5 <= my_rom(6751); 
 data6 <= my_rom(8106); 
 data7 <= my_rom(9461); 
 data8 <= my_rom(10816); 
 data9 <= my_rom(12171); 
 data10 <= my_rom(13526);
when "10100110100" => 
 data1 <= my_rom(1332); 
 data2 <= my_rom(2687); 
 data3 <= my_rom(4042); 
 data4 <= my_rom(5397); 
 data5 <= my_rom(6752); 
 data6 <= my_rom(8107); 
 data7 <= my_rom(9462); 
 data8 <= my_rom(10817); 
 data9 <= my_rom(12172); 
 data10 <= my_rom(13527);
when "10100110101" => 
 data1 <= my_rom(1333); 
 data2 <= my_rom(2688); 
 data3 <= my_rom(4043); 
 data4 <= my_rom(5398); 
 data5 <= my_rom(6753); 
 data6 <= my_rom(8108); 
 data7 <= my_rom(9463); 
 data8 <= my_rom(10818); 
 data9 <= my_rom(12173); 
 data10 <= my_rom(13528);
when "10100110110" => 
 data1 <= my_rom(1334); 
 data2 <= my_rom(2689); 
 data3 <= my_rom(4044); 
 data4 <= my_rom(5399); 
 data5 <= my_rom(6754); 
 data6 <= my_rom(8109); 
 data7 <= my_rom(9464); 
 data8 <= my_rom(10819); 
 data9 <= my_rom(12174); 
 data10 <= my_rom(13529);
when "10100110111" => 
 data1 <= my_rom(1335); 
 data2 <= my_rom(2690); 
 data3 <= my_rom(4045); 
 data4 <= my_rom(5400); 
 data5 <= my_rom(6755); 
 data6 <= my_rom(8110); 
 data7 <= my_rom(9465); 
 data8 <= my_rom(10820); 
 data9 <= my_rom(12175); 
 data10 <= my_rom(13530);
when "10100111000" => 
 data1 <= my_rom(1336); 
 data2 <= my_rom(2691); 
 data3 <= my_rom(4046); 
 data4 <= my_rom(5401); 
 data5 <= my_rom(6756); 
 data6 <= my_rom(8111); 
 data7 <= my_rom(9466); 
 data8 <= my_rom(10821); 
 data9 <= my_rom(12176); 
 data10 <= my_rom(13531);
when "10100111001" => 
 data1 <= my_rom(1337); 
 data2 <= my_rom(2692); 
 data3 <= my_rom(4047); 
 data4 <= my_rom(5402); 
 data5 <= my_rom(6757); 
 data6 <= my_rom(8112); 
 data7 <= my_rom(9467); 
 data8 <= my_rom(10822); 
 data9 <= my_rom(12177); 
 data10 <= my_rom(13532);
when "10100111010" => 
 data1 <= my_rom(1338); 
 data2 <= my_rom(2693); 
 data3 <= my_rom(4048); 
 data4 <= my_rom(5403); 
 data5 <= my_rom(6758); 
 data6 <= my_rom(8113); 
 data7 <= my_rom(9468); 
 data8 <= my_rom(10823); 
 data9 <= my_rom(12178); 
 data10 <= my_rom(13533);
when "10100111011" => 
 data1 <= my_rom(1339); 
 data2 <= my_rom(2694); 
 data3 <= my_rom(4049); 
 data4 <= my_rom(5404); 
 data5 <= my_rom(6759); 
 data6 <= my_rom(8114); 
 data7 <= my_rom(9469); 
 data8 <= my_rom(10824); 
 data9 <= my_rom(12179); 
 data10 <= my_rom(13534);
when "10100111100" => 
 data1 <= my_rom(1340); 
 data2 <= my_rom(2695); 
 data3 <= my_rom(4050); 
 data4 <= my_rom(5405); 
 data5 <= my_rom(6760); 
 data6 <= my_rom(8115); 
 data7 <= my_rom(9470); 
 data8 <= my_rom(10825); 
 data9 <= my_rom(12180); 
 data10 <= my_rom(13535);
when "10100111101" => 
 data1 <= my_rom(1341); 
 data2 <= my_rom(2696); 
 data3 <= my_rom(4051); 
 data4 <= my_rom(5406); 
 data5 <= my_rom(6761); 
 data6 <= my_rom(8116); 
 data7 <= my_rom(9471); 
 data8 <= my_rom(10826); 
 data9 <= my_rom(12181); 
 data10 <= my_rom(13536);
when "10100111110" => 
 data1 <= my_rom(1342); 
 data2 <= my_rom(2697); 
 data3 <= my_rom(4052); 
 data4 <= my_rom(5407); 
 data5 <= my_rom(6762); 
 data6 <= my_rom(8117); 
 data7 <= my_rom(9472); 
 data8 <= my_rom(10827); 
 data9 <= my_rom(12182); 
 data10 <= my_rom(13537);
when "10100111111" => 
 data1 <= my_rom(1343); 
 data2 <= my_rom(2698); 
 data3 <= my_rom(4053); 
 data4 <= my_rom(5408); 
 data5 <= my_rom(6763); 
 data6 <= my_rom(8118); 
 data7 <= my_rom(9473); 
 data8 <= my_rom(10828); 
 data9 <= my_rom(12183); 
 data10 <= my_rom(13538);
when "10101000000" => 
 data1 <= my_rom(1344); 
 data2 <= my_rom(2699); 
 data3 <= my_rom(4054); 
 data4 <= my_rom(5409); 
 data5 <= my_rom(6764); 
 data6 <= my_rom(8119); 
 data7 <= my_rom(9474); 
 data8 <= my_rom(10829); 
 data9 <= my_rom(12184); 
 data10 <= my_rom(13539);
when "10101000001" => 
 data1 <= my_rom(1345); 
 data2 <= my_rom(2700); 
 data3 <= my_rom(4055); 
 data4 <= my_rom(5410); 
 data5 <= my_rom(6765); 
 data6 <= my_rom(8120); 
 data7 <= my_rom(9475); 
 data8 <= my_rom(10830); 
 data9 <= my_rom(12185); 
 data10 <= my_rom(13540);
when "10101000010" => 
 data1 <= my_rom(1346); 
 data2 <= my_rom(2701); 
 data3 <= my_rom(4056); 
 data4 <= my_rom(5411); 
 data5 <= my_rom(6766); 
 data6 <= my_rom(8121); 
 data7 <= my_rom(9476); 
 data8 <= my_rom(10831); 
 data9 <= my_rom(12186); 
 data10 <= my_rom(13541);
when "10101000011" => 
 data1 <= my_rom(1347); 
 data2 <= my_rom(2702); 
 data3 <= my_rom(4057); 
 data4 <= my_rom(5412); 
 data5 <= my_rom(6767); 
 data6 <= my_rom(8122); 
 data7 <= my_rom(9477); 
 data8 <= my_rom(10832); 
 data9 <= my_rom(12187); 
 data10 <= my_rom(13542);
when "10101000100" => 
 data1 <= my_rom(1348); 
 data2 <= my_rom(2703); 
 data3 <= my_rom(4058); 
 data4 <= my_rom(5413); 
 data5 <= my_rom(6768); 
 data6 <= my_rom(8123); 
 data7 <= my_rom(9478); 
 data8 <= my_rom(10833); 
 data9 <= my_rom(12188); 
 data10 <= my_rom(13543);
when "10101000101" => 
 data1 <= my_rom(1349); 
 data2 <= my_rom(2704); 
 data3 <= my_rom(4059); 
 data4 <= my_rom(5414); 
 data5 <= my_rom(6769); 
 data6 <= my_rom(8124); 
 data7 <= my_rom(9479); 
 data8 <= my_rom(10834); 
 data9 <= my_rom(12189); 
 data10 <= my_rom(13544);
when "10101000110" => 
 data1 <= my_rom(1350); 
 data2 <= my_rom(2705); 
 data3 <= my_rom(4060); 
 data4 <= my_rom(5415); 
 data5 <= my_rom(6770); 
 data6 <= my_rom(8125); 
 data7 <= my_rom(9480); 
 data8 <= my_rom(10835); 
 data9 <= my_rom(12190); 
 data10 <= my_rom(13545);
when "10101000111" => 
 data1 <= my_rom(1351); 
 data2 <= my_rom(2706); 
 data3 <= my_rom(4061); 
 data4 <= my_rom(5416); 
 data5 <= my_rom(6771); 
 data6 <= my_rom(8126); 
 data7 <= my_rom(9481); 
 data8 <= my_rom(10836); 
 data9 <= my_rom(12191); 
 data10 <= my_rom(13546);
when "10101001000" => 
 data1 <= my_rom(1352); 
 data2 <= my_rom(2707); 
 data3 <= my_rom(4062); 
 data4 <= my_rom(5417); 
 data5 <= my_rom(6772); 
 data6 <= my_rom(8127); 
 data7 <= my_rom(9482); 
 data8 <= my_rom(10837); 
 data9 <= my_rom(12192); 
 data10 <= my_rom(13547);
when "10101001001" => 
 data1 <= my_rom(1353); 
 data2 <= my_rom(2708); 
 data3 <= my_rom(4063); 
 data4 <= my_rom(5418); 
 data5 <= my_rom(6773); 
 data6 <= my_rom(8128); 
 data7 <= my_rom(9483); 
 data8 <= my_rom(10838); 
 data9 <= my_rom(12193); 
 data10 <= my_rom(13548);
when others => 
 data1 <= my_rom(1354); 
 data2 <= my_rom(2709); 
 data3 <= my_rom(4064); 
 data4 <= my_rom(5419); 
 data5 <= my_rom(6774); 
 data6 <= my_rom(8129); 
 data7 <= my_rom(9484); 
 data8 <= my_rom(10839); 
 data9 <= my_rom(12194); 
 data10 <= my_rom(13549);
    end case;
end process;
end behavioral;